// rom.v
// to be included from the top module at the compile

initial
begin
    mem['h0000]=8'hC0; mem['h0001]=8'h44; mem['h0002]=8'hB6; mem['h0003]=8'h08;
    mem['h0004]=8'hFF; mem['h0005]=8'hFF; mem['h0006]=8'hFF; mem['h0007]=8'hFF;
    mem['h0008]=8'hFF; mem['h0009]=8'hFF; mem['h000A]=8'hFF; mem['h000B]=8'hFF;
    mem['h000C]=8'hFF; mem['h000D]=8'hFF; mem['h000E]=8'hFF; mem['h000F]=8'hFF;
    mem['h0010]=8'hFF; mem['h0011]=8'hFF; mem['h0012]=8'hFF; mem['h0013]=8'hFF;
    mem['h0014]=8'hFF; mem['h0015]=8'hFF; mem['h0016]=8'hFF; mem['h0017]=8'hFF;
    mem['h0018]=8'hFF; mem['h0019]=8'hFF; mem['h001A]=8'hFF; mem['h001B]=8'hFF;
    mem['h001C]=8'hFF; mem['h001D]=8'hFF; mem['h001E]=8'hFF; mem['h001F]=8'hFF;
    mem['h0020]=8'hFF; mem['h0021]=8'hFF; mem['h0022]=8'hFF; mem['h0023]=8'hFF;
    mem['h0024]=8'hFF; mem['h0025]=8'hFF; mem['h0026]=8'hFF; mem['h0027]=8'hFF;
    mem['h0028]=8'hFF; mem['h0029]=8'hFF; mem['h002A]=8'hFF; mem['h002B]=8'hFF;
    mem['h002C]=8'hFF; mem['h002D]=8'hFF; mem['h002E]=8'hFF; mem['h002F]=8'hFF;
    mem['h0030]=8'hFF; mem['h0031]=8'hFF; mem['h0032]=8'hFF; mem['h0033]=8'hFF;
    mem['h0034]=8'hFF; mem['h0035]=8'hFF; mem['h0036]=8'hFF; mem['h0037]=8'hFF;
    mem['h0038]=8'hFF; mem['h0039]=8'hFF; mem['h003A]=8'hFF; mem['h003B]=8'hFF;
    mem['h003C]=8'hFF; mem['h003D]=8'hFF; mem['h003E]=8'hFF; mem['h003F]=8'hFF;
    mem['h0040]=8'h44; mem['h0041]=8'hB6; mem['h0042]=8'h08; mem['h0043]=8'h41;
    mem['h0044]=8'h1A; mem['h0045]=8'h40; mem['h0046]=8'h43; mem['h0047]=8'h00;
    mem['h0048]=8'h43; mem['h0049]=8'h61; mem['h004A]=8'h34; mem['h004B]=8'h80;
    mem['h004C]=8'h07; mem['h004D]=8'h00; mem['h004E]=8'hC8; mem['h004F]=8'h24;
    mem['h0050]=8'h7F; mem['h0051]=8'h3C; mem['h0052]=8'h0D; mem['h0053]=8'h68;
    mem['h0054]=8'h65; mem['h0055]=8'h00; mem['h0056]=8'h3C; mem['h0057]=8'h0A;
    mem['h0058]=8'h68; mem['h0059]=8'h65; mem['h005A]=8'h00; mem['h005B]=8'h3C;
    mem['h005C]=8'h7F; mem['h005D]=8'h68; mem['h005E]=8'h68; mem['h005F]=8'h00;
    mem['h0060]=8'h3C; mem['h0061]=8'h20; mem['h0062]=8'h60; mem['h0063]=8'h68;
    mem['h0064]=8'h00; mem['h0065]=8'h61; mem['h0066]=8'hC1; mem['h0067]=8'h07;
    mem['h0068]=8'h06; mem['h0069]=8'h3C; mem['h006A]=8'h61; mem['h006B]=8'hC1;
    mem['h006C]=8'h1A; mem['h006D]=8'h1A; mem['h006E]=8'h1A; mem['h006F]=8'h1A;
    mem['h0070]=8'h24; mem['h0071]=8'h0F; mem['h0072]=8'h04; mem['h0073]=8'h30;
    mem['h0074]=8'h3C; mem['h0075]=8'h3A; mem['h0076]=8'h60; mem['h0077]=8'h7B;
    mem['h0078]=8'h00; mem['h0079]=8'h04; mem['h007A]=8'h07; mem['h007B]=8'h61;
    mem['h007C]=8'hC1; mem['h007D]=8'h24; mem['h007E]=8'h0F; mem['h007F]=8'h04;
    mem['h0080]=8'h30; mem['h0081]=8'h3C; mem['h0082]=8'h3A; mem['h0083]=8'h60;
    mem['h0084]=8'h88; mem['h0085]=8'h00; mem['h0086]=8'h04; mem['h0087]=8'h07;
    mem['h0088]=8'h61; mem['h0089]=8'h06; mem['h008A]=8'h3E; mem['h008B]=8'h61;
    mem['h008C]=8'hC1; mem['h008D]=8'h07; mem['h008E]=8'hFF; mem['h008F]=8'hFF;
    mem['h0090]=8'hFF; mem['h0091]=8'hFF; mem['h0092]=8'hFF; mem['h0093]=8'hFF;
    mem['h0094]=8'hFF; mem['h0095]=8'hFF; mem['h0096]=8'hFF; mem['h0097]=8'hFF;
    mem['h0098]=8'hFF; mem['h0099]=8'hFF; mem['h009A]=8'hFF; mem['h009B]=8'hFF;
    mem['h009C]=8'hFF; mem['h009D]=8'hFF; mem['h009E]=8'hFF; mem['h009F]=8'hFF;
    mem['h00A0]=8'hFF; mem['h00A1]=8'hFF; mem['h00A2]=8'hFF; mem['h00A3]=8'hFF;
    mem['h00A4]=8'hFF; mem['h00A5]=8'hFF; mem['h00A6]=8'hFF; mem['h00A7]=8'hFF;
    mem['h00A8]=8'hFF; mem['h00A9]=8'hFF; mem['h00AA]=8'hFF; mem['h00AB]=8'hFF;
    mem['h00AC]=8'hFF; mem['h00AD]=8'hFF; mem['h00AE]=8'hFF; mem['h00AF]=8'hFF;
    mem['h00B0]=8'hFF; mem['h00B1]=8'hFF; mem['h00B2]=8'hFF; mem['h00B3]=8'hFF;
    mem['h00B4]=8'hFF; mem['h00B5]=8'hFF; mem['h00B6]=8'hFF; mem['h00B7]=8'hFF;
    mem['h00B8]=8'hFF; mem['h00B9]=8'hFF; mem['h00BA]=8'hFF; mem['h00BB]=8'hFF;
    mem['h00BC]=8'hFF; mem['h00BD]=8'hFF; mem['h00BE]=8'hFF; mem['h00BF]=8'hFF;
    mem['h00C0]=8'hFF; mem['h00C1]=8'hFF; mem['h00C2]=8'hFF; mem['h00C3]=8'hFF;
    mem['h00C4]=8'hFF; mem['h00C5]=8'hFF; mem['h00C6]=8'hFF; mem['h00C7]=8'hFF;
    mem['h00C8]=8'hFF; mem['h00C9]=8'hFF; mem['h00CA]=8'hFF; mem['h00CB]=8'hFF;
    mem['h00CC]=8'hFF; mem['h00CD]=8'hFF; mem['h00CE]=8'hFF; mem['h00CF]=8'hFF;
    mem['h00D0]=8'hFF; mem['h00D1]=8'hFF; mem['h00D2]=8'hFF; mem['h00D3]=8'hFF;
    mem['h00D4]=8'hFF; mem['h00D5]=8'hFF; mem['h00D6]=8'hFF; mem['h00D7]=8'hFF;
    mem['h00D8]=8'hFF; mem['h00D9]=8'hFF; mem['h00DA]=8'hFF; mem['h00DB]=8'hFF;
    mem['h00DC]=8'hFF; mem['h00DD]=8'hFF; mem['h00DE]=8'hFF; mem['h00DF]=8'hFF;
    mem['h00E0]=8'hFF; mem['h00E1]=8'hFF; mem['h00E2]=8'hFF; mem['h00E3]=8'hFF;
    mem['h00E4]=8'hFF; mem['h00E5]=8'hFF; mem['h00E6]=8'hFF; mem['h00E7]=8'hFF;
    mem['h00E8]=8'hFF; mem['h00E9]=8'hFF; mem['h00EA]=8'hFF; mem['h00EB]=8'hFF;
    mem['h00EC]=8'hFF; mem['h00ED]=8'hFF; mem['h00EE]=8'hFF; mem['h00EF]=8'hFF;
    mem['h00F0]=8'hFF; mem['h00F1]=8'hFF; mem['h00F2]=8'hFF; mem['h00F3]=8'hFF;
    mem['h00F4]=8'hFF; mem['h00F5]=8'hFF; mem['h00F6]=8'hFF; mem['h00F7]=8'hFF;
    mem['h00F8]=8'hFF; mem['h00F9]=8'hFF; mem['h00FA]=8'hFF; mem['h00FB]=8'hFF;
    mem['h00FC]=8'hFF; mem['h00FD]=8'hFF; mem['h00FE]=8'hFF; mem['h00FF]=8'hFF;
    mem['h0100]=8'hFF; mem['h0101]=8'hFF; mem['h0102]=8'hFF; mem['h0103]=8'hFF;
    mem['h0104]=8'h00; mem['h0105]=8'h00; mem['h0106]=8'h40; mem['h0107]=8'h01;
    mem['h0108]=8'hFF; mem['h0109]=8'hFF; mem['h010A]=8'hFF; mem['h010B]=8'h00;
    mem['h010C]=8'h00; mem['h010D]=8'h00; mem['h010E]=8'h00; mem['h010F]=8'h00;
    mem['h0110]=8'hFF; mem['h0111]=8'hFF; mem['h0112]=8'hFF; mem['h0113]=8'hFF;
    mem['h0114]=8'h00; mem['h0115]=8'h00; mem['h0116]=8'hC0; mem['h0117]=8'h01;
    mem['h0118]=8'h00; mem['h0119]=8'h00; mem['h011A]=8'h00; mem['h011B]=8'h00;
    mem['h011C]=8'h00; mem['h011D]=8'h00; mem['h011E]=8'h00; mem['h011F]=8'h00;
    mem['h0120]=8'h00; mem['h0121]=8'h00; mem['h0122]=8'h00; mem['h0123]=8'h00;
    mem['h0124]=8'h00; mem['h0125]=8'h00; mem['h0126]=8'h00; mem['h0127]=8'h00;
    mem['h0128]=8'h01; mem['h0129]=8'h50; mem['h012A]=8'h72; mem['h012B]=8'h02;
    mem['h012C]=8'hFF; mem['h012D]=8'hFF; mem['h012E]=8'hFF; mem['h012F]=8'hFF;
    mem['h0130]=8'h03; mem['h0131]=8'h68; mem['h0132]=8'h6F; mem['h0133]=8'h0C;
    mem['h0134]=8'h00; mem['h0135]=8'h00; mem['h0136]=8'h00; mem['h0137]=8'h00;
    mem['h0138]=8'h00; mem['h0139]=8'h00; mem['h013A]=8'h00; mem['h013B]=8'h00;
    mem['h013C]=8'h00; mem['h013D]=8'h00; mem['h013E]=8'h00; mem['h013F]=8'h00;
    mem['h0140]=8'h00; mem['h0141]=8'h00; mem['h0142]=8'h00; mem['h0143]=8'h00;
    mem['h0144]=8'h00; mem['h0145]=8'h00; mem['h0146]=8'h00; mem['h0147]=8'h00;
    mem['h0148]=8'h00; mem['h0149]=8'hFF; mem['h014A]=8'hFF; mem['h014B]=8'hFF;
    mem['h014C]=8'hFF; mem['h014D]=8'hFF; mem['h014E]=8'hFF; mem['h014F]=8'hFF;
    mem['h0150]=8'h00; mem['h0151]=8'h00; mem['h0152]=8'h00; mem['h0153]=8'h00;
    mem['h0154]=8'h00; mem['h0155]=8'h00; mem['h0156]=8'h00; mem['h0157]=8'h00;
    mem['h0158]=8'h00; mem['h0159]=8'h00; mem['h015A]=8'h00; mem['h015B]=8'h00;
    mem['h015C]=8'h00; mem['h015D]=8'h00; mem['h015E]=8'h00; mem['h015F]=8'h00;
    mem['h0160]=8'h00; mem['h0161]=8'h00; mem['h0162]=8'h00; mem['h0163]=8'h00;
    mem['h0164]=8'h00; mem['h0165]=8'h00; mem['h0166]=8'h00; mem['h0167]=8'h00;
    mem['h0168]=8'h00; mem['h0169]=8'h00; mem['h016A]=8'h00; mem['h016B]=8'h00;
    mem['h016C]=8'h00; mem['h016D]=8'h00; mem['h016E]=8'h00; mem['h016F]=8'h00;
    mem['h0170]=8'h00; mem['h0171]=8'h00; mem['h0172]=8'h00; mem['h0173]=8'h00;
    mem['h0174]=8'h00; mem['h0175]=8'h00; mem['h0176]=8'h00; mem['h0177]=8'h00;
    mem['h0178]=8'hFF; mem['h0179]=8'hFF; mem['h017A]=8'hFF; mem['h017B]=8'hFF;
    mem['h017C]=8'hFF; mem['h017D]=8'hFF; mem['h017E]=8'hFF; mem['h017F]=8'hFF;
    mem['h0180]=8'h00; mem['h0181]=8'h00; mem['h0182]=8'h00; mem['h0183]=8'h00;
    mem['h0184]=8'hFF; mem['h0185]=8'hFF; mem['h0186]=8'hFF; mem['h0187]=8'hFF;
    mem['h0188]=8'h00; mem['h0189]=8'h00; mem['h018A]=8'h50; mem['h018B]=8'h04;
    mem['h018C]=8'h67; mem['h018D]=8'h66; mem['h018E]=8'h66; mem['h018F]=8'hFD;
    mem['h0190]=8'h00; mem['h0191]=8'hFF; mem['h0192]=8'hFF; mem['h0193]=8'hFF;
    mem['h0194]=8'hFF; mem['h0195]=8'hFF; mem['h0196]=8'hFF; mem['h0197]=8'h00;
    mem['h0198]=8'h00; mem['h0199]=8'hFF; mem['h019A]=8'hFF; mem['h019B]=8'hFF;
    mem['h019C]=8'hFF; mem['h019D]=8'hFF; mem['h019E]=8'hFF; mem['h019F]=8'hFF;
    mem['h01A0]=8'hFF; mem['h01A1]=8'hFF; mem['h01A2]=8'hFF; mem['h01A3]=8'hFF;
    mem['h01A4]=8'hFF; mem['h01A5]=8'hFF; mem['h01A6]=8'hFF; mem['h01A7]=8'hFF;
    mem['h01A8]=8'hFF; mem['h01A9]=8'hFF; mem['h01AA]=8'hFF; mem['h01AB]=8'hFF;
    mem['h01AC]=8'hFF; mem['h01AD]=8'hFF; mem['h01AE]=8'hFF; mem['h01AF]=8'hFF;
    mem['h01B0]=8'hFF; mem['h01B1]=8'hFF; mem['h01B2]=8'hFF; mem['h01B3]=8'hFF;
    mem['h01B4]=8'hFF; mem['h01B5]=8'hFF; mem['h01B6]=8'hFF; mem['h01B7]=8'hFF;
    mem['h01B8]=8'hFF; mem['h01B9]=8'hFF; mem['h01BA]=8'h04; mem['h01BB]=8'hD3;
    mem['h01BC]=8'hC1; mem['h01BD]=8'hD6; mem['h01BE]=8'hC5; mem['h01BF]=8'h04;
    mem['h01C0]=8'hCC; mem['h01C1]=8'hCF; mem['h01C2]=8'hC1; mem['h01C3]=8'hC4;
    mem['h01C4]=8'h00; mem['h01C5]=8'h00; mem['h01C6]=8'h00; mem['h01C7]=8'h00;
    mem['h01C8]=8'h00; mem['h01C9]=8'h00; mem['h01CA]=8'h00; mem['h01CB]=8'h00;
    mem['h01CC]=8'h00; mem['h01CD]=8'h00; mem['h01CE]=8'h00; mem['h01CF]=8'h00;
    mem['h01D0]=8'h04; mem['h01D1]=8'hD4; mem['h01D2]=8'hC8; mem['h01D3]=8'hC5;
    mem['h01D4]=8'hCE; mem['h01D5]=8'h02; mem['h01D6]=8'hD4; mem['h01D7]=8'hCF;
    mem['h01D8]=8'h04; mem['h01D9]=8'hD3; mem['h01DA]=8'hD4; mem['h01DB]=8'hC5;
    mem['h01DC]=8'hD0; mem['h01DD]=8'h04; mem['h01DE]=8'hCC; mem['h01DF]=8'hC9;
    mem['h01E0]=8'hD3; mem['h01E1]=8'hD4; mem['h01E2]=8'h03; mem['h01E3]=8'hD2;
    mem['h01E4]=8'hD5; mem['h01E5]=8'hCE; mem['h01E6]=8'h03; mem['h01E7]=8'hD3;
    mem['h01E8]=8'hC3; mem['h01E9]=8'hD2; mem['h01EA]=8'h0B; mem['h01EB]=8'h8D;
    mem['h01EC]=8'h8D; mem['h01ED]=8'h8A; mem['h01EE]=8'hD2; mem['h01EF]=8'hC5;
    mem['h01F0]=8'hC1; mem['h01F1]=8'hC4; mem['h01F2]=8'hD9; mem['h01F3]=8'h8D;
    mem['h01F4]=8'h8A; mem['h01F5]=8'h8A; mem['h01F6]=8'h09; mem['h01F7]=8'hA0;
    mem['h01F8]=8'hC1; mem['h01F9]=8'hD4; mem['h01FA]=8'hA0; mem['h01FB]=8'hCC;
    mem['h01FC]=8'hC9; mem['h01FD]=8'hCE; mem['h01FE]=8'hC5; mem['h01FF]=8'hA0;
    mem['h0200]=8'h46; mem['h0201]=8'hAD; mem['h0202]=8'h02; mem['h0203]=8'h36;
    mem['h0204]=8'hE0; mem['h0205]=8'h2E; mem['h0206]=8'h16; mem['h0207]=8'h3E;
    mem['h0208]=8'h00; mem['h0209]=8'h36; mem['h020A]=8'h81; mem['h020B]=8'h3E;
    mem['h020C]=8'h01; mem['h020D]=8'h36; mem['h020E]=8'h81; mem['h020F]=8'h46;
    mem['h0210]=8'hA0; mem['h0211]=8'h02; mem['h0212]=8'h68; mem['h0213]=8'h24;
    mem['h0214]=8'h02; mem['h0215]=8'h3C; mem['h0216]=8'hB0; mem['h0217]=8'h70;
    mem['h0218]=8'h31; mem['h0219]=8'h02; mem['h021A]=8'h3C; mem['h021B]=8'hBA;
    mem['h021C]=8'h50; mem['h021D]=8'h31; mem['h021E]=8'h02; mem['h021F]=8'h36;
    mem['h0220]=8'hE0; mem['h0221]=8'h46; mem['h0222]=8'hCC; mem['h0223]=8'h02;
    mem['h0224]=8'h36; mem['h0225]=8'h81; mem['h0226]=8'h46; mem['h0227]=8'h03;
    mem['h0228]=8'h03; mem['h0229]=8'h48; mem['h022A]=8'h0D; mem['h022B]=8'h02;
    mem['h022C]=8'h36; mem['h022D]=8'h83; mem['h022E]=8'h3E; mem['h022F]=8'h00;
    mem['h0230]=8'h07; mem['h0231]=8'h36; mem['h0232]=8'h81; mem['h0233]=8'hCF;
    mem['h0234]=8'h36; mem['h0235]=8'h82; mem['h0236]=8'hF9; mem['h0237]=8'h36;
    mem['h0238]=8'h82; mem['h0239]=8'h46; mem['h023A]=8'hA0; mem['h023B]=8'h02;
    mem['h023C]=8'h68; mem['h023D]=8'h79; mem['h023E]=8'h02; mem['h023F]=8'h3C;
    mem['h0240]=8'hBD; mem['h0241]=8'h68; mem['h0242]=8'h88; mem['h0243]=8'h02;
    mem['h0244]=8'h3C; mem['h0245]=8'hA8; mem['h0246]=8'h68; mem['h0247]=8'h8D;
    mem['h0248]=8'h02; mem['h0249]=8'h46; mem['h024A]=8'hC8; mem['h024B]=8'h02;
    mem['h024C]=8'h36; mem['h024D]=8'h83; mem['h024E]=8'h3E; mem['h024F]=8'h01;
    mem['h0250]=8'h2E; mem['h0251]=8'h17; mem['h0252]=8'h36; mem['h0253]=8'h00;
    mem['h0254]=8'h1E; mem['h0255]=8'h16; mem['h0256]=8'h26; mem['h0257]=8'h50;
    mem['h0258]=8'h46; mem['h0259]=8'hDA; mem['h025A]=8'h02; mem['h025B]=8'h2B;
    mem['h025C]=8'h46; mem['h025D]=8'hEE; mem['h025E]=8'h12; mem['h025F]=8'h30;
    mem['h0260]=8'hC7; mem['h0261]=8'h24; mem['h0262]=8'hC0; mem['h0263]=8'h48;
    mem['h0264]=8'h5F; mem['h0265]=8'h02; mem['h0266]=8'h46; mem['h0267]=8'hEE;
    mem['h0268]=8'h12; mem['h0269]=8'h36; mem['h026A]=8'h83; mem['h026B]=8'h2E;
    mem['h026C]=8'h16; mem['h026D]=8'hCF; mem['h026E]=8'h08; mem['h026F]=8'hF9;
    mem['h0270]=8'h46; mem['h0271]=8'hEE; mem['h0272]=8'h12; mem['h0273]=8'hC1;
    mem['h0274]=8'h3C; mem['h0275]=8'h0D; mem['h0276]=8'h48; mem['h0277]=8'h54;
    mem['h0278]=8'h02; mem['h0279]=8'h36; mem['h027A]=8'h82; mem['h027B]=8'h2E;
    mem['h027C]=8'h16; mem['h027D]=8'h46; mem['h027E]=8'h03; mem['h027F]=8'h03;
    mem['h0280]=8'h48; mem['h0281]=8'h37; mem['h0282]=8'h02; mem['h0283]=8'h36;
    mem['h0284]=8'h83; mem['h0285]=8'h3E; mem['h0286]=8'hFF; mem['h0287]=8'h07;
    mem['h0288]=8'h36; mem['h0289]=8'h83; mem['h028A]=8'h3E; mem['h028B]=8'h0D;
    mem['h028C]=8'h07; mem['h028D]=8'h36; mem['h028E]=8'h83; mem['h028F]=8'h3E;
    mem['h0290]=8'h0E; mem['h0291]=8'h07; mem['h0292]=8'h06; mem['h0293]=8'hC2;
    mem['h0294]=8'h16; mem['h0295]=8'hC7; mem['h0296]=8'h46; mem['h0297]=8'h82;
    mem['h0298]=8'h03; mem['h0299]=8'hC2; mem['h029A]=8'h46; mem['h029B]=8'h82;
    mem['h029C]=8'h03; mem['h029D]=8'h44; mem['h029E]=8'hD2; mem['h029F]=8'h0A;
    mem['h02A0]=8'hC7; mem['h02A1]=8'h3C; mem['h02A2]=8'h50; mem['h02A3]=8'h50;
    mem['h02A4]=8'h92; mem['h02A5]=8'h02; mem['h02A6]=8'hF0; mem['h02A7]=8'h2E;
    mem['h02A8]=8'h16; mem['h02A9]=8'hC7; mem['h02AA]=8'h3C; mem['h02AB]=8'hA0;
    mem['h02AC]=8'h07; mem['h02AD]=8'h36; mem['h02AE]=8'h50; mem['h02AF]=8'h2E;
    mem['h02B0]=8'h16; mem['h02B1]=8'h3E; mem['h02B2]=8'h00; mem['h02B3]=8'h07;
    mem['h02B4]=8'h3C; mem['h02B5]=8'hC1; mem['h02B6]=8'h70; mem['h02B7]=8'hBE;
    mem['h02B8]=8'h02; mem['h02B9]=8'h3C; mem['h02BA]=8'hDB; mem['h02BB]=8'h70;
    mem['h02BC]=8'hC8; mem['h02BD]=8'h02; mem['h02BE]=8'h3C; mem['h02BF]=8'hB0;
    mem['h02C0]=8'h70; mem['h02C1]=8'hD7; mem['h02C2]=8'h02; mem['h02C3]=8'h3C;
    mem['h02C4]=8'hBA; mem['h02C5]=8'h50; mem['h02C6]=8'hD7; mem['h02C7]=8'h02;
    mem['h02C8]=8'h36; mem['h02C9]=8'h50; mem['h02CA]=8'h2E; mem['h02CB]=8'h16;
    mem['h02CC]=8'hD7; mem['h02CD]=8'h10; mem['h02CE]=8'hFA; mem['h02CF]=8'hC8;
    mem['h02D0]=8'h46; mem['h02D1]=8'h1E; mem['h02D2]=8'h13; mem['h02D3]=8'hF9;
    mem['h02D4]=8'h06; mem['h02D5]=8'h00; mem['h02D6]=8'h07; mem['h02D7]=8'h44;
    mem['h02D8]=8'h6A; mem['h02D9]=8'h09; mem['h02DA]=8'hC7; mem['h02DB]=8'h46;
    mem['h02DC]=8'hEE; mem['h02DD]=8'h12; mem['h02DE]=8'hCF; mem['h02DF]=8'hB9;
    mem['h02E0]=8'h0B; mem['h02E1]=8'h46; mem['h02E2]=8'hEE; mem['h02E3]=8'h12;
    mem['h02E4]=8'h46; mem['h02E5]=8'hFF; mem['h02E6]=8'h02; mem['h02E7]=8'hC7;
    mem['h02E8]=8'h46; mem['h02E9]=8'hEE; mem['h02EA]=8'h12; mem['h02EB]=8'h46;
    mem['h02EC]=8'hFF; mem['h02ED]=8'h02; mem['h02EE]=8'hBF; mem['h02EF]=8'h0B;
    mem['h02F0]=8'h46; mem['h02F1]=8'hEE; mem['h02F2]=8'h12; mem['h02F3]=8'h09;
    mem['h02F4]=8'h48; mem['h02F5]=8'hE4; mem['h02F6]=8'h02; mem['h02F7]=8'h07;
    mem['h02F8]=8'hC7; mem['h02F9]=8'h46; mem['h02FA]=8'hEE; mem['h02FB]=8'h12;
    mem['h02FC]=8'h44; mem['h02FD]=8'hEE; mem['h02FE]=8'h02; mem['h02FF]=8'h30;
    mem['h0300]=8'h0B; mem['h0301]=8'h28; mem['h0302]=8'h07; mem['h0303]=8'hCF;
    mem['h0304]=8'h08; mem['h0305]=8'hF9; mem['h0306]=8'h36; mem['h0307]=8'h00;
    mem['h0308]=8'hC7; mem['h0309]=8'h09; mem['h030A]=8'hB9; mem['h030B]=8'h07;
    mem['h030C]=8'h16; mem['h030D]=8'h00; mem['h030E]=8'h46; mem['h030F]=8'h91;
    mem['h0310]=8'h03; mem['h0311]=8'h3C; mem['h0312]=8'hFF; mem['h0313]=8'h48;
    mem['h0314]=8'h25; mem['h0315]=8'h03; mem['h0316]=8'h06; mem['h0317]=8'hDC;
    mem['h0318]=8'h46; mem['h0319]=8'h82; mem['h031A]=8'h03; mem['h031B]=8'h11;
    mem['h031C]=8'h70; mem['h031D]=8'h0C; mem['h031E]=8'h03; mem['h031F]=8'h46;
    mem['h0320]=8'h74; mem['h0321]=8'h03; mem['h0322]=8'h44; mem['h0323]=8'h0E;
    mem['h0324]=8'h03; mem['h0325]=8'h3C; mem['h0326]=8'h83; mem['h0327]=8'h68;
    mem['h0328]=8'hCB; mem['h0329]=8'h0A; mem['h032A]=8'h3C; mem['h032B]=8'h8D;
    mem['h032C]=8'h68; mem['h032D]=8'h42; mem['h032E]=8'h03; mem['h032F]=8'h3C;
    mem['h0330]=8'h8A; mem['h0331]=8'h68; mem['h0332]=8'h0E; mem['h0333]=8'h03;
    mem['h0334]=8'h46; mem['h0335]=8'hFF; mem['h0336]=8'h02; mem['h0337]=8'h10;
    mem['h0338]=8'hF8; mem['h0339]=8'hC2; mem['h033A]=8'h3C; mem['h033B]=8'h50;
    mem['h033C]=8'h50; mem['h033D]=8'h92; mem['h033E]=8'h02; mem['h033F]=8'h44;
    mem['h0340]=8'h0E; mem['h0341]=8'h03; mem['h0342]=8'hCA; mem['h0343]=8'h46;
    mem['h0344]=8'h4B; mem['h0345]=8'h03; mem['h0346]=8'hFA; mem['h0347]=8'h46;
    mem['h0348]=8'h61; mem['h0349]=8'h03; mem['h034A]=8'h07; mem['h034B]=8'hC6;
    mem['h034C]=8'h91; mem['h034D]=8'hF0; mem['h034E]=8'h03; mem['h034F]=8'h29;
    mem['h0350]=8'h07; mem['h0351]=8'hD7; mem['h0352]=8'hC7; mem['h0353]=8'hA0;
    mem['h0354]=8'h2B; mem['h0355]=8'h46; mem['h0356]=8'hFF; mem['h0357]=8'h02;
    mem['h0358]=8'hC7; mem['h0359]=8'h46; mem['h035A]=8'h82; mem['h035B]=8'h03;
    mem['h035C]=8'h11; mem['h035D]=8'h48; mem['h035E]=8'h55; mem['h035F]=8'h03;
    mem['h0360]=8'h07; mem['h0361]=8'h06; mem['h0362]=8'h8D; mem['h0363]=8'h46;
    mem['h0364]=8'h82; mem['h0365]=8'h03; mem['h0366]=8'h06; mem['h0367]=8'h8A;
    mem['h0368]=8'h46; mem['h0369]=8'h82; mem['h036A]=8'h03; mem['h036B]=8'h36;
    mem['h036C]=8'h23; mem['h036D]=8'h2E; mem['h036E]=8'h01; mem['h036F]=8'h3E;
    mem['h0370]=8'h01; mem['h0371]=8'hEB; mem['h0372]=8'hF4; mem['h0373]=8'h07;
    mem['h0374]=8'h31; mem['h0375]=8'h30; mem['h0376]=8'h48; mem['h0377]=8'h7A;
    mem['h0378]=8'h03; mem['h0379]=8'h29; mem['h037A]=8'h31; mem['h037B]=8'h07;
    mem['h037C]=8'hC6; mem['h037D]=8'h81; mem['h037E]=8'hF0; mem['h037F]=8'h03;
    mem['h0380]=8'h28; mem['h0381]=8'h07; mem['h0382]=8'hDD; mem['h0383]=8'hE6;
    mem['h0384]=8'h36; mem['h0385]=8'h23; mem['h0386]=8'h2E; mem['h0387]=8'h01;
    mem['h0388]=8'hCF; mem['h0389]=8'h08; mem['h038A]=8'hF9; mem['h038B]=8'h46;
    mem['h038C]=8'h4E; mem['h038D]=8'h00; mem['h038E]=8'hEB; mem['h038F]=8'hF4;
    mem['h0390]=8'h07; mem['h0391]=8'h44; mem['h0392]=8'h43; mem['h0393]=8'h00;
    mem['h0394]=8'h36; mem['h0395]=8'h97; mem['h0396]=8'h2E; mem['h0397]=8'h01;
    mem['h0398]=8'h3E; mem['h0399]=8'h94; mem['h039A]=8'h30; mem['h039B]=8'h2E;
    mem['h039C]=8'h16; mem['h039D]=8'h3E; mem['h039E]=8'h00; mem['h039F]=8'h46;
    mem['h03A0]=8'hAD; mem['h03A1]=8'h02; mem['h03A2]=8'h36; mem['h03A3]=8'h88;
    mem['h03A4]=8'h3E; mem['h03A5]=8'h00; mem['h03A6]=8'h36; mem['h03A7]=8'hBE;
    mem['h03A8]=8'hCF; mem['h03A9]=8'h36; mem['h03AA]=8'h80; mem['h03AB]=8'hF9;
    mem['h03AC]=8'h36; mem['h03AD]=8'h80; mem['h03AE]=8'h46; mem['h03AF]=8'hA0;
    mem['h03B0]=8'h02; mem['h03B1]=8'h68; mem['h03B2]=8'hC1; mem['h03B3]=8'h04;
    mem['h03B4]=8'h3C; mem['h03B5]=8'hAB; mem['h03B6]=8'h48; mem['h03B7]=8'hC0;
    mem['h03B8]=8'h03; mem['h03B9]=8'h36; mem['h03BA]=8'h7E; mem['h03BB]=8'h3E;
    mem['h03BC]=8'h01; mem['h03BD]=8'h44; mem['h03BE]=8'hE9; mem['h03BF]=8'h03;
    mem['h03C0]=8'h3C; mem['h03C1]=8'hAD; mem['h03C2]=8'h48; mem['h03C3]=8'hEF;
    mem['h03C4]=8'h03; mem['h03C5]=8'h36; mem['h03C6]=8'h50; mem['h03C7]=8'hC7;
    mem['h03C8]=8'hA0; mem['h03C9]=8'h48; mem['h03CA]=8'hE5; mem['h03CB]=8'h03;
    mem['h03CC]=8'h36; mem['h03CD]=8'h7E; mem['h03CE]=8'hC7; mem['h03CF]=8'h3C;
    mem['h03D0]=8'h07; mem['h03D1]=8'h68; mem['h03D2]=8'hE5; mem['h03D3]=8'h03;
    mem['h03D4]=8'h3C; mem['h03D5]=8'h03; mem['h03D6]=8'h68; mem['h03D7]=8'h6A;
    mem['h03D8]=8'h09; mem['h03D9]=8'h3C; mem['h03DA]=8'h05; mem['h03DB]=8'h68;
    mem['h03DC]=8'h6A; mem['h03DD]=8'h09; mem['h03DE]=8'h36; mem['h03DF]=8'h50;
    mem['h03E0]=8'h3E; mem['h03E1]=8'h01; mem['h03E2]=8'h30; mem['h03E3]=8'h3E;
    mem['h03E4]=8'hB0; mem['h03E5]=8'h36; mem['h03E6]=8'h7E; mem['h03E7]=8'h3E;
    mem['h03E8]=8'h02; mem['h03E9]=8'h46; mem['h03EA]=8'hD4; mem['h03EB]=8'h04;
    mem['h03EC]=8'h44; mem['h03ED]=8'hC1; mem['h03EE]=8'h04; mem['h03EF]=8'h3C;
    mem['h03F0]=8'hAA; mem['h03F1]=8'h48; mem['h03F2]=8'hFB; mem['h03F3]=8'h03;
    mem['h03F4]=8'h36; mem['h03F5]=8'h7E; mem['h03F6]=8'h3E; mem['h03F7]=8'h03;
    mem['h03F8]=8'h44; mem['h03F9]=8'hE9; mem['h03FA]=8'h03; mem['h03FB]=8'h3C;
    mem['h03FC]=8'hAF; mem['h03FD]=8'h48; mem['h03FE]=8'h07; mem['h03FF]=8'h04;
    mem['h0400]=8'h36; mem['h0401]=8'h7E; mem['h0402]=8'h3E; mem['h0403]=8'h04;
    mem['h0404]=8'h44; mem['h0405]=8'hE9; mem['h0406]=8'h03; mem['h0407]=8'h3C;
    mem['h0408]=8'hA8; mem['h0409]=8'h48; mem['h040A]=8'h1B; mem['h040B]=8'h04;
    mem['h040C]=8'h36; mem['h040D]=8'h98; mem['h040E]=8'hCF; mem['h040F]=8'h08;
    mem['h0410]=8'hF9; mem['h0411]=8'h46; mem['h0412]=8'h40; mem['h0413]=8'h07;
    mem['h0414]=8'h36; mem['h0415]=8'h7E; mem['h0416]=8'h3E; mem['h0417]=8'h06;
    mem['h0418]=8'h44; mem['h0419]=8'hE9; mem['h041A]=8'h03; mem['h041B]=8'h3C;
    mem['h041C]=8'hA9; mem['h041D]=8'h48; mem['h041E]=8'h34; mem['h041F]=8'h04;
    mem['h0420]=8'h36; mem['h0421]=8'h7E; mem['h0422]=8'h3E; mem['h0423]=8'h07;
    mem['h0424]=8'h46; mem['h0425]=8'hD4; mem['h0426]=8'h04; mem['h0427]=8'h46;
    mem['h0428]=8'h03; mem['h0429]=8'h07; mem['h042A]=8'h36; mem['h042B]=8'h98;
    mem['h042C]=8'h2E; mem['h042D]=8'h16; mem['h042E]=8'hCF; mem['h042F]=8'h09;
    mem['h0430]=8'hF9; mem['h0431]=8'h44; mem['h0432]=8'hC1; mem['h0433]=8'h04;
    mem['h0434]=8'h3C; mem['h0435]=8'hDE; mem['h0436]=8'h48; mem['h0437]=8'h40;
    mem['h0438]=8'h04; mem['h0439]=8'h36; mem['h043A]=8'h7E; mem['h043B]=8'h3E;
    mem['h043C]=8'h05; mem['h043D]=8'h44; mem['h043E]=8'hE9; mem['h043F]=8'h03;
    mem['h0440]=8'h3C; mem['h0441]=8'hBC; mem['h0442]=8'h48; mem['h0443]=8'h63;
    mem['h0444]=8'h04; mem['h0445]=8'h36; mem['h0446]=8'h80; mem['h0447]=8'hCF;
    mem['h0448]=8'h08; mem['h0449]=8'hF9; mem['h044A]=8'h46; mem['h044B]=8'hA0;
    mem['h044C]=8'h02; mem['h044D]=8'h3C; mem['h044E]=8'hBD; mem['h044F]=8'h68;
    mem['h0450]=8'hA9; mem['h0451]=8'h04; mem['h0452]=8'h3C; mem['h0453]=8'hBE;
    mem['h0454]=8'h68; mem['h0455]=8'hB7; mem['h0456]=8'h04; mem['h0457]=8'h36;
    mem['h0458]=8'h80; mem['h0459]=8'hCF; mem['h045A]=8'h09; mem['h045B]=8'hF9;
    mem['h045C]=8'h36; mem['h045D]=8'h7E; mem['h045E]=8'h3E; mem['h045F]=8'h09;
    mem['h0460]=8'h44; mem['h0461]=8'hE9; mem['h0462]=8'h03; mem['h0463]=8'h3C;
    mem['h0464]=8'hBD; mem['h0465]=8'h48; mem['h0466]=8'h86; mem['h0467]=8'h04;
    mem['h0468]=8'h36; mem['h0469]=8'h80; mem['h046A]=8'hCF; mem['h046B]=8'h08;
    mem['h046C]=8'hF9; mem['h046D]=8'h46; mem['h046E]=8'hA0; mem['h046F]=8'h02;
    mem['h0470]=8'h3C; mem['h0471]=8'hBC; mem['h0472]=8'h68; mem['h0473]=8'hA9;
    mem['h0474]=8'h04; mem['h0475]=8'h3C; mem['h0476]=8'hBE; mem['h0477]=8'h68;
    mem['h0478]=8'hB0; mem['h0479]=8'h04; mem['h047A]=8'h36; mem['h047B]=8'h80;
    mem['h047C]=8'hCF; mem['h047D]=8'h09; mem['h047E]=8'hF9; mem['h047F]=8'h36;
    mem['h0480]=8'h7E; mem['h0481]=8'h3E; mem['h0482]=8'h0A; mem['h0483]=8'h44;
    mem['h0484]=8'hE9; mem['h0485]=8'h03; mem['h0486]=8'h3C; mem['h0487]=8'hBE;
    mem['h0488]=8'h48; mem['h0489]=8'hBE; mem['h048A]=8'h04; mem['h048B]=8'h36;
    mem['h048C]=8'h80; mem['h048D]=8'hCF; mem['h048E]=8'h08; mem['h048F]=8'hF9;
    mem['h0490]=8'h46; mem['h0491]=8'hA0; mem['h0492]=8'h02; mem['h0493]=8'h3C;
    mem['h0494]=8'hBC; mem['h0495]=8'h68; mem['h0496]=8'hB7; mem['h0497]=8'h04;
    mem['h0498]=8'h3C; mem['h0499]=8'hBD; mem['h049A]=8'h68; mem['h049B]=8'hB0;
    mem['h049C]=8'h04; mem['h049D]=8'h36; mem['h049E]=8'h80; mem['h049F]=8'hCF;
    mem['h04A0]=8'h09; mem['h04A1]=8'hF9; mem['h04A2]=8'h36; mem['h04A3]=8'h7E;
    mem['h04A4]=8'h3E; mem['h04A5]=8'h0B; mem['h04A6]=8'h44; mem['h04A7]=8'hE9;
    mem['h04A8]=8'h03; mem['h04A9]=8'h36; mem['h04AA]=8'h7E; mem['h04AB]=8'h3E;
    mem['h04AC]=8'h0C; mem['h04AD]=8'h44; mem['h04AE]=8'hE9; mem['h04AF]=8'h03;
    mem['h04B0]=8'h36; mem['h04B1]=8'h7E; mem['h04B2]=8'h3E; mem['h04B3]=8'h0D;
    mem['h04B4]=8'h44; mem['h04B5]=8'hE9; mem['h04B6]=8'h03; mem['h04B7]=8'h36;
    mem['h04B8]=8'h7E; mem['h04B9]=8'h3E; mem['h04BA]=8'h0E; mem['h04BB]=8'h44;
    mem['h04BC]=8'hE9; mem['h04BD]=8'h03; mem['h04BE]=8'h46; mem['h04BF]=8'hC8;
    mem['h04C0]=8'h02; mem['h04C1]=8'h36; mem['h04C2]=8'h80; mem['h04C3]=8'h2E;
    mem['h04C4]=8'h16; mem['h04C5]=8'hCF; mem['h04C6]=8'h08; mem['h04C7]=8'hF9;
    mem['h04C8]=8'h36; mem['h04C9]=8'hBF; mem['h04CA]=8'hC7; mem['h04CB]=8'h09;
    mem['h04CC]=8'hB9; mem['h04CD]=8'h48; mem['h04CE]=8'hAC; mem['h04CF]=8'h03;
    mem['h04D0]=8'h44; mem['h04D1]=8'hC0; mem['h04D2]=8'h19; mem['h04D3]=8'h00;
    mem['h04D4]=8'h36; mem['h04D5]=8'h50; mem['h04D6]=8'h2E; mem['h04D7]=8'h16;
    mem['h04D8]=8'hC7; mem['h04D9]=8'hA0; mem['h04DA]=8'h68; mem['h04DB]=8'h99;
    mem['h04DC]=8'h05; mem['h04DD]=8'h30; mem['h04DE]=8'hC7; mem['h04DF]=8'h3C;
    mem['h04E0]=8'hAE; mem['h04E1]=8'h68; mem['h04E2]=8'hEE; mem['h04E3]=8'h04;
    mem['h04E4]=8'h3C; mem['h04E5]=8'hB0; mem['h04E6]=8'h70; mem['h04E7]=8'h1B;
    mem['h04E8]=8'h05; mem['h04E9]=8'h3C; mem['h04EA]=8'hBA; mem['h04EB]=8'h50;
    mem['h04EC]=8'h1B; mem['h04ED]=8'h05; mem['h04EE]=8'h31; mem['h04EF]=8'hC7;
    mem['h04F0]=8'h3C; mem['h04F1]=8'h01; mem['h04F2]=8'h68; mem['h04F3]=8'h05;
    mem['h04F4]=8'h05; mem['h04F5]=8'h86; mem['h04F6]=8'hF0; mem['h04F7]=8'hC7;
    mem['h04F8]=8'h3C; mem['h04F9]=8'hC5; mem['h04FA]=8'h48; mem['h04FB]=8'h05;
    mem['h04FC]=8'h05; mem['h04FD]=8'h36; mem['h04FE]=8'h80; mem['h04FF]=8'h46;
    mem['h0500]=8'hA0; mem['h0501]=8'h02; mem['h0502]=8'h44; mem['h0503]=8'hC8;
    mem['h0504]=8'h02; mem['h0505]=8'h36; mem['h0506]=8'h97; mem['h0507]=8'h2E;
    mem['h0508]=8'h01; mem['h0509]=8'hC7; mem['h050A]=8'h04; mem['h050B]=8'h04;
    mem['h050C]=8'hF8; mem['h050D]=8'hF0; mem['h050E]=8'h46; mem['h050F]=8'hAD;
    mem['h0510]=8'h12; mem['h0511]=8'h36; mem['h0512]=8'h50; mem['h0513]=8'h2E;
    mem['h0514]=8'h16; mem['h0515]=8'h46; mem['h0516]=8'h24; mem['h0517]=8'h13;
    mem['h0518]=8'h44; mem['h0519]=8'h99; mem['h051A]=8'h05; mem['h051B]=8'h36;
    mem['h051C]=8'hF8; mem['h051D]=8'h2E; mem['h051E]=8'h16; mem['h051F]=8'h3E;
    mem['h0520]=8'h00; mem['h0521]=8'h36; mem['h0522]=8'h50; mem['h0523]=8'h1E;
    mem['h0524]=8'h17; mem['h0525]=8'h26; mem['h0526]=8'h88; mem['h0527]=8'hC7;
    mem['h0528]=8'h3C; mem['h0529]=8'h01; mem['h052A]=8'h48; mem['h052B]=8'h31;
    mem['h052C]=8'h05; mem['h052D]=8'h36; mem['h052E]=8'h52; mem['h052F]=8'h3E;
    mem['h0530]=8'h00; mem['h0531]=8'h36; mem['h0532]=8'h51; mem['h0533]=8'h2E;
    mem['h0534]=8'h16; mem['h0535]=8'h46; mem['h0536]=8'hEE; mem['h0537]=8'h12;
    mem['h0538]=8'hC7; mem['h0539]=8'h30; mem['h053A]=8'hCF; mem['h053B]=8'h30;
    mem['h053C]=8'h46; mem['h053D]=8'hEE; mem['h053E]=8'h12; mem['h053F]=8'hBF;
    mem['h0540]=8'h48; mem['h0541]=8'h49; mem['h0542]=8'h05; mem['h0543]=8'h30;
    mem['h0544]=8'hC1; mem['h0545]=8'hBF; mem['h0546]=8'h68; mem['h0547]=8'h81;
    mem['h0548]=8'h05; mem['h0549]=8'h46; mem['h054A]=8'hAE; mem['h054B]=8'h06;
    mem['h054C]=8'h36; mem['h054D]=8'hF8; mem['h054E]=8'h2E; mem['h054F]=8'h16;
    mem['h0550]=8'hCF; mem['h0551]=8'h08; mem['h0552]=8'hF9; mem['h0553]=8'h36;
    mem['h0554]=8'h3F; mem['h0555]=8'h2E; mem['h0556]=8'h17; mem['h0557]=8'hC1;
    mem['h0558]=8'hBF; mem['h0559]=8'h48; mem['h055A]=8'h31; mem['h055B]=8'h05;
    mem['h055C]=8'h36; mem['h055D]=8'h3F; mem['h055E]=8'h2E; mem['h055F]=8'h17;
    mem['h0560]=8'hCF; mem['h0561]=8'h08; mem['h0562]=8'hF9; mem['h0563]=8'hC1;
    mem['h0564]=8'h3C; mem['h0565]=8'h15; mem['h0566]=8'h50; mem['h0567]=8'h92;
    mem['h0568]=8'h02; mem['h0569]=8'h36; mem['h056A]=8'h51; mem['h056B]=8'h2E;
    mem['h056C]=8'h16; mem['h056D]=8'h0E; mem['h056E]=8'h02; mem['h056F]=8'h46;
    mem['h0570]=8'h0B; mem['h0571]=8'h11; mem['h0572]=8'hF4; mem['h0573]=8'hEB;
    mem['h0574]=8'hA8; mem['h0575]=8'hF8; mem['h0576]=8'h30; mem['h0577]=8'hF8;
    mem['h0578]=8'h30; mem['h0579]=8'hF8; mem['h057A]=8'h30; mem['h057B]=8'hF8;
    mem['h057C]=8'hC6; mem['h057D]=8'h14; mem['h057E]=8'h04; mem['h057F]=8'hE0;
    mem['h0580]=8'hDD; mem['h0581]=8'h46; mem['h0582]=8'hCF; mem['h0583]=8'h12;
    mem['h0584]=8'h36; mem['h0585]=8'h97; mem['h0586]=8'h2E; mem['h0587]=8'h01;
    mem['h0588]=8'hC7; mem['h0589]=8'h04; mem['h058A]=8'h04; mem['h058B]=8'hF8;
    mem['h058C]=8'hF0; mem['h058D]=8'h46; mem['h058E]=8'hAD; mem['h058F]=8'h12;
    mem['h0590]=8'h46; mem['h0591]=8'hDF; mem['h0592]=8'h12; mem['h0593]=8'h46;
    mem['h0594]=8'hEE; mem['h0595]=8'h12; mem['h0596]=8'h46; mem['h0597]=8'hA4;
    mem['h0598]=8'h12; mem['h0599]=8'h46; mem['h059A]=8'hAD; mem['h059B]=8'h02;
    mem['h059C]=8'h36; mem['h059D]=8'h7E; mem['h059E]=8'hC7; mem['h059F]=8'h3C;
    mem['h05A0]=8'h07; mem['h05A1]=8'h68; mem['h05A2]=8'hDA; mem['h05A3]=8'h05;
    mem['h05A4]=8'h04; mem['h05A5]=8'hA0; mem['h05A6]=8'hF0; mem['h05A7]=8'hCF;
    mem['h05A8]=8'h36; mem['h05A9]=8'h88; mem['h05AA]=8'hD7; mem['h05AB]=8'h46;
    mem['h05AC]=8'h1E; mem['h05AD]=8'h13; mem['h05AE]=8'hC7; mem['h05AF]=8'h04;
    mem['h05B0]=8'hAF; mem['h05B1]=8'hF0; mem['h05B2]=8'hC1; mem['h05B3]=8'hBF;
    mem['h05B4]=8'h68; mem['h05B5]=8'hC7; mem['h05B6]=8'h05; mem['h05B7]=8'h70;
    mem['h05B8]=8'hC7; mem['h05B9]=8'h05; mem['h05BA]=8'h36; mem['h05BB]=8'h7E;
    mem['h05BC]=8'hCF; mem['h05BD]=8'h36; mem['h05BE]=8'h88; mem['h05BF]=8'hD7;
    mem['h05C0]=8'h10; mem['h05C1]=8'hFA; mem['h05C2]=8'h46; mem['h05C3]=8'h1E;
    mem['h05C4]=8'h13; mem['h05C5]=8'hF9; mem['h05C6]=8'h07; mem['h05C7]=8'h36;
    mem['h05C8]=8'h88; mem['h05C9]=8'hC7; mem['h05CA]=8'h86; mem['h05CB]=8'hF0;
    mem['h05CC]=8'hC7; mem['h05CD]=8'hA0; mem['h05CE]=8'h2B; mem['h05CF]=8'h36;
    mem['h05D0]=8'h88; mem['h05D1]=8'hD7; mem['h05D2]=8'h11; mem['h05D3]=8'hFA;
    mem['h05D4]=8'h46; mem['h05D5]=8'hF4; mem['h05D6]=8'h05; mem['h05D7]=8'h44;
    mem['h05D8]=8'h99; mem['h05D9]=8'h05; mem['h05DA]=8'h36; mem['h05DB]=8'h88;
    mem['h05DC]=8'h2E; mem['h05DD]=8'h16; mem['h05DE]=8'hC7; mem['h05DF]=8'h86;
    mem['h05E0]=8'hF0; mem['h05E1]=8'hC7; mem['h05E2]=8'hA0; mem['h05E3]=8'h68;
    mem['h05E4]=8'h44; mem['h05E5]=8'h06; mem['h05E6]=8'h36; mem['h05E7]=8'h88;
    mem['h05E8]=8'hD7; mem['h05E9]=8'h11; mem['h05EA]=8'hFA; mem['h05EB]=8'h3C;
    mem['h05EC]=8'h06; mem['h05ED]=8'h2B; mem['h05EE]=8'h46; mem['h05EF]=8'hF4;
    mem['h05F0]=8'h05; mem['h05F1]=8'h44; mem['h05F2]=8'hDA; mem['h05F3]=8'h05;
    mem['h05F4]=8'h36; mem['h05F5]=8'hF9; mem['h05F6]=8'h2E; mem['h05F7]=8'h16;
    mem['h05F8]=8'hF8; mem['h05F9]=8'h36; mem['h05FA]=8'h97; mem['h05FB]=8'h2E;
    mem['h05FC]=8'h01; mem['h05FD]=8'hC7; mem['h05FE]=8'hF0; mem['h05FF]=8'h46;
    mem['h0600]=8'hB6; mem['h0601]=8'h12; mem['h0602]=8'h36; mem['h0603]=8'h97;
    mem['h0604]=8'hC7; mem['h0605]=8'h14; mem['h0606]=8'h04; mem['h0607]=8'hF8;
    mem['h0608]=8'h36; mem['h0609]=8'hF9; mem['h060A]=8'h2E; mem['h060B]=8'h16;
    mem['h060C]=8'hC7; mem['h060D]=8'h3C; mem['h060E]=8'h01; mem['h060F]=8'h68;
    mem['h0610]=8'h89; mem['h0611]=8'h10; mem['h0612]=8'h3C; mem['h0613]=8'h02;
    mem['h0614]=8'h68; mem['h0615]=8'h1A; mem['h0616]=8'h11; mem['h0617]=8'h3C;
    mem['h0618]=8'h03; mem['h0619]=8'h68; mem['h061A]=8'h26; mem['h061B]=8'h11;
    mem['h061C]=8'h3C; mem['h061D]=8'h04; mem['h061E]=8'h68; mem['h061F]=8'hD2;
    mem['h0620]=8'h11; mem['h0621]=8'h3C; mem['h0622]=8'h05; mem['h0623]=8'h68;
    mem['h0624]=8'hB3; mem['h0625]=8'h06; mem['h0626]=8'h3C; mem['h0627]=8'h09;
    mem['h0628]=8'h68; mem['h0629]=8'h51; mem['h062A]=8'h06; mem['h062B]=8'h3C;
    mem['h062C]=8'h0A; mem['h062D]=8'h68; mem['h062E]=8'h5E; mem['h062F]=8'h06;
    mem['h0630]=8'h3C; mem['h0631]=8'h0B; mem['h0632]=8'h68; mem['h0633]=8'h6B;
    mem['h0634]=8'h06; mem['h0635]=8'h3C; mem['h0636]=8'h0C; mem['h0637]=8'h68;
    mem['h0638]=8'h7B; mem['h0639]=8'h06; mem['h063A]=8'h3C; mem['h063B]=8'h0D;
    mem['h063C]=8'h68; mem['h063D]=8'h8B; mem['h063E]=8'h06; mem['h063F]=8'h3C;
    mem['h0640]=8'h0E; mem['h0641]=8'h68; mem['h0642]=8'h98; mem['h0643]=8'h06;
    mem['h0644]=8'h36; mem['h0645]=8'h98; mem['h0646]=8'h2E; mem['h0647]=8'h16;
    mem['h0648]=8'h3E; mem['h0649]=8'h00; mem['h064A]=8'h06; mem['h064B]=8'hC9;
    mem['h064C]=8'h16; mem['h064D]=8'hA8; mem['h064E]=8'h44; mem['h064F]=8'h96;
    mem['h0650]=8'h02; mem['h0651]=8'h46; mem['h0652]=8'h1A; mem['h0653]=8'h11;
    mem['h0654]=8'h36; mem['h0655]=8'h56; mem['h0656]=8'hC7; mem['h0657]=8'hA0;
    mem['h0658]=8'h70; mem['h0659]=8'hA2; mem['h065A]=8'h06; mem['h065B]=8'h44;
    mem['h065C]=8'hA7; mem['h065D]=8'h06; mem['h065E]=8'h46; mem['h065F]=8'h1A;
    mem['h0660]=8'h11; mem['h0661]=8'h36; mem['h0662]=8'h56; mem['h0663]=8'hC7;
    mem['h0664]=8'hA0; mem['h0665]=8'h68; mem['h0666]=8'hA2; mem['h0667]=8'h06;
    mem['h0668]=8'h44; mem['h0669]=8'hA7; mem['h066A]=8'h06; mem['h066B]=8'h46;
    mem['h066C]=8'h1A; mem['h066D]=8'h11; mem['h066E]=8'h36; mem['h066F]=8'h56;
    mem['h0670]=8'hC7; mem['h0671]=8'hA0; mem['h0672]=8'h68; mem['h0673]=8'hA7;
    mem['h0674]=8'h06; mem['h0675]=8'h50; mem['h0676]=8'hA2; mem['h0677]=8'h06;
    mem['h0678]=8'h44; mem['h0679]=8'hA7; mem['h067A]=8'h06; mem['h067B]=8'h46;
    mem['h067C]=8'h1A; mem['h067D]=8'h11; mem['h067E]=8'h36; mem['h067F]=8'h56;
    mem['h0680]=8'hC7; mem['h0681]=8'hA0; mem['h0682]=8'h68; mem['h0683]=8'hA2;
    mem['h0684]=8'h06; mem['h0685]=8'h70; mem['h0686]=8'hA2; mem['h0687]=8'h06;
    mem['h0688]=8'h44; mem['h0689]=8'hA7; mem['h068A]=8'h06; mem['h068B]=8'h46;
    mem['h068C]=8'h1A; mem['h068D]=8'h11; mem['h068E]=8'h36; mem['h068F]=8'h56;
    mem['h0690]=8'hC7; mem['h0691]=8'hA0; mem['h0692]=8'h50; mem['h0693]=8'hA2;
    mem['h0694]=8'h06; mem['h0695]=8'h44; mem['h0696]=8'hA7; mem['h0697]=8'h06;
    mem['h0698]=8'h46; mem['h0699]=8'h1A; mem['h069A]=8'h11; mem['h069B]=8'h36;
    mem['h069C]=8'h56; mem['h069D]=8'hC7; mem['h069E]=8'hA0; mem['h069F]=8'h68;
    mem['h06A0]=8'hA7; mem['h06A1]=8'h06; mem['h06A2]=8'h36; mem['h06A3]=8'h04;
    mem['h06A4]=8'h44; mem['h06A5]=8'hA4; mem['h06A6]=8'h12; mem['h06A7]=8'h36;
    mem['h06A8]=8'h57; mem['h06A9]=8'h3E; mem['h06AA]=8'h00; mem['h06AB]=8'h44;
    mem['h06AC]=8'h29; mem['h06AD]=8'h10; mem['h06AE]=8'hC4; mem['h06AF]=8'h04;
    mem['h06B0]=8'h04; mem['h06B1]=8'hE0; mem['h06B2]=8'h07; mem['h06B3]=8'h36;
    mem['h06B4]=8'h56; mem['h06B5]=8'h2E; mem['h06B6]=8'h01; mem['h06B7]=8'hC7;
    mem['h06B8]=8'h36; mem['h06B9]=8'h03; mem['h06BA]=8'hF8; mem['h06BB]=8'hA0;
    mem['h06BC]=8'h68; mem['h06BD]=8'hA2; mem['h06BE]=8'h06; mem['h06BF]=8'h72;
    mem['h06C0]=8'h82; mem['h06C1]=8'h10; mem['h06C2]=8'h46; mem['h06C3]=8'h00;
    mem['h06C4]=8'h10; mem['h06C5]=8'h36; mem['h06C6]=8'h54; mem['h06C7]=8'hCF;
    mem['h06C8]=8'h36; mem['h06C9]=8'h0B; mem['h06CA]=8'hF9; mem['h06CB]=8'h36;
    mem['h06CC]=8'h5C; mem['h06CD]=8'h26; mem['h06CE]=8'h0C; mem['h06CF]=8'h2E;
    mem['h06D0]=8'h01; mem['h06D1]=8'hDD; mem['h06D2]=8'h0E; mem['h06D3]=8'h04;
    mem['h06D4]=8'h46; mem['h06D5]=8'h0B; mem['h06D6]=8'h11; mem['h06D7]=8'h46;
    mem['h06D8]=8'hA2; mem['h06D9]=8'h06; mem['h06DA]=8'h36; mem['h06DB]=8'h03;
    mem['h06DC]=8'hC7; mem['h06DD]=8'hA0; mem['h06DE]=8'h70; mem['h06DF]=8'hF2;
    mem['h06E0]=8'h06; mem['h06E1]=8'h36; mem['h06E2]=8'h0C; mem['h06E3]=8'h46;
    mem['h06E4]=8'hBF; mem['h06E5]=8'h12; mem['h06E6]=8'h46; mem['h06E7]=8'h26;
    mem['h06E8]=8'h11; mem['h06E9]=8'h36; mem['h06EA]=8'h0B; mem['h06EB]=8'hCF;
    mem['h06EC]=8'h09; mem['h06ED]=8'hF9; mem['h06EE]=8'h48; mem['h06EF]=8'hE1;
    mem['h06F0]=8'h06; mem['h06F1]=8'h07; mem['h06F2]=8'h36; mem['h06F3]=8'h0C;
    mem['h06F4]=8'h46; mem['h06F5]=8'hBF; mem['h06F6]=8'h12; mem['h06F7]=8'h46;
    mem['h06F8]=8'hD2; mem['h06F9]=8'h11; mem['h06FA]=8'h36; mem['h06FB]=8'h0B;
    mem['h06FC]=8'hCF; mem['h06FD]=8'h09; mem['h06FE]=8'hF9; mem['h06FF]=8'h48;
    mem['h0700]=8'hF2; mem['h0701]=8'h06; mem['h0702]=8'h07; mem['h0703]=8'h36;
    mem['h0704]=8'h98; mem['h0705]=8'h2E; mem['h0706]=8'h16; mem['h0707]=8'hC7;
    mem['h0708]=8'h86; mem['h0709]=8'hF0; mem['h070A]=8'hC7; mem['h070B]=8'h3E;
    mem['h070C]=8'h00; mem['h070D]=8'h36; mem['h070E]=8'h83; mem['h070F]=8'h2E;
    mem['h0710]=8'h17; mem['h0711]=8'hF8; mem['h0712]=8'hA0; mem['h0713]=8'h2B;
    mem['h0714]=8'h70; mem['h0715]=8'h00; mem['h0716]=8'h2D; mem['h0717]=8'h3C;
    mem['h0718]=8'h01; mem['h0719]=8'h68; mem['h071A]=8'hA3; mem['h071B]=8'h07;
    mem['h071C]=8'h3C; mem['h071D]=8'h02; mem['h071E]=8'h68; mem['h071F]=8'hF0;
    mem['h0720]=8'h07; mem['h0721]=8'h3C; mem['h0722]=8'h03; mem['h0723]=8'h68;
    mem['h0724]=8'hE6; mem['h0725]=8'h07; mem['h0726]=8'h3C; mem['h0727]=8'h04;
    mem['h0728]=8'h68; mem['h0729]=8'h00; mem['h072A]=8'h1A; mem['h072B]=8'h3C;
    mem['h072C]=8'h05; mem['h072D]=8'h68; mem['h072E]=8'h0F; mem['h072F]=8'h08;
    mem['h0730]=8'h3C; mem['h0731]=8'h06; mem['h0732]=8'h68; mem['h0733]=8'hA0;
    mem['h0734]=8'h1A; mem['h0735]=8'h3C; mem['h0736]=8'h07; mem['h0737]=8'h68;
    mem['h0738]=8'hFF; mem['h0739]=8'h07; mem['h073A]=8'h3C; mem['h073B]=8'h08;
    mem['h073C]=8'h68; mem['h073D]=8'h4D; mem['h073E]=8'h00; mem['h073F]=8'h00;
    mem['h0740]=8'h36; mem['h0741]=8'h50; mem['h0742]=8'h2E; mem['h0743]=8'h16;
    mem['h0744]=8'hC7; mem['h0745]=8'hA0; mem['h0746]=8'h2B; mem['h0747]=8'h36;
    mem['h0748]=8'h82; mem['h0749]=8'h2E; mem['h074A]=8'h17; mem['h074B]=8'h3E;
    mem['h074C]=8'h00; mem['h074D]=8'h36; mem['h074E]=8'h82; mem['h074F]=8'h2E;
    mem['h0750]=8'h17; mem['h0751]=8'hCF; mem['h0752]=8'h08; mem['h0753]=8'hF9;
    mem['h0754]=8'h16; mem['h0755]=8'h02; mem['h0756]=8'h36; mem['h0757]=8'hBC;
    mem['h0758]=8'h2E; mem['h0759]=8'h16; mem['h075A]=8'h46; mem['h075B]=8'h98;
    mem['h075C]=8'h07; mem['h075D]=8'h1E; mem['h075E]=8'h16; mem['h075F]=8'h26;
    mem['h0760]=8'h50; mem['h0761]=8'h46; mem['h0762]=8'hDA; mem['h0763]=8'h02;
    mem['h0764]=8'h68; mem['h0765]=8'h87; mem['h0766]=8'h07; mem['h0767]=8'h36;
    mem['h0768]=8'h82; mem['h0769]=8'h2E; mem['h076A]=8'h17; mem['h076B]=8'hC7;
    mem['h076C]=8'h3C; mem['h076D]=8'h08; mem['h076E]=8'h48; mem['h076F]=8'h4D;
    mem['h0770]=8'h07; mem['h0771]=8'h36; mem['h0772]=8'h82; mem['h0773]=8'h2E;
    mem['h0774]=8'h17; mem['h0775]=8'h3E; mem['h0776]=8'h00; mem['h0777]=8'h44;
    mem['h0778]=8'h2C; mem['h0779]=8'h2D; mem['h077A]=8'h36; mem['h077B]=8'h98;
    mem['h077C]=8'h2E; mem['h077D]=8'h16; mem['h077E]=8'h3E; mem['h077F]=8'h00;
    mem['h0780]=8'h06; mem['h0781]=8'hC6; mem['h0782]=8'h16; mem['h0783]=8'hC1;
    mem['h0784]=8'h44; mem['h0785]=8'h96; mem['h0786]=8'h02; mem['h0787]=8'h36;
    mem['h0788]=8'h82; mem['h0789]=8'h2E; mem['h078A]=8'h17; mem['h078B]=8'hCF;
    mem['h078C]=8'h36; mem['h078D]=8'h98; mem['h078E]=8'h2E; mem['h078F]=8'h16;
    mem['h0790]=8'hD7; mem['h0791]=8'h46; mem['h0792]=8'h1E; mem['h0793]=8'h13;
    mem['h0794]=8'hF9; mem['h0795]=8'h44; mem['h0796]=8'hAD; mem['h0797]=8'h02;
    mem['h0798]=8'hC1; mem['h0799]=8'h02; mem['h079A]=8'h11; mem['h079B]=8'h48;
    mem['h079C]=8'h99; mem['h079D]=8'h07; mem['h079E]=8'h86; mem['h079F]=8'hF0;
    mem['h07A0]=8'h03; mem['h07A1]=8'h28; mem['h07A2]=8'h07; mem['h07A3]=8'h36;
    mem['h07A4]=8'h56; mem['h07A5]=8'h2E; mem['h07A6]=8'h01; mem['h07A7]=8'hC7;
    mem['h07A8]=8'hA0; mem['h07A9]=8'h50; mem['h07AA]=8'hD7; mem['h07AB]=8'h07;
    mem['h07AC]=8'h36; mem['h07AD]=8'h0C; mem['h07AE]=8'h46; mem['h07AF]=8'hAD;
    mem['h07B0]=8'h12; mem['h07B1]=8'h46; mem['h07B2]=8'h00; mem['h07B3]=8'h10;
    mem['h07B4]=8'h36; mem['h07B5]=8'h53; mem['h07B6]=8'h3E; mem['h07B7]=8'h00;
    mem['h07B8]=8'h46; mem['h07B9]=8'h34; mem['h07BA]=8'h10; mem['h07BB]=8'h36;
    mem['h07BC]=8'h0C; mem['h07BD]=8'h46; mem['h07BE]=8'hB6; mem['h07BF]=8'h12;
    mem['h07C0]=8'h46; mem['h07C1]=8'h1A; mem['h07C2]=8'h11; mem['h07C3]=8'h36;
    mem['h07C4]=8'h56; mem['h07C5]=8'hC7; mem['h07C6]=8'hA0; mem['h07C7]=8'h68;
    mem['h07C8]=8'hE1; mem['h07C9]=8'h07; mem['h07CA]=8'h36; mem['h07CB]=8'h0C;
    mem['h07CC]=8'h46; mem['h07CD]=8'hA4; mem['h07CE]=8'h12; mem['h07CF]=8'h36;
    mem['h07D0]=8'h14; mem['h07D1]=8'h46; mem['h07D2]=8'hBF; mem['h07D3]=8'h12;
    mem['h07D4]=8'h46; mem['h07D5]=8'h89; mem['h07D6]=8'h10; mem['h07D7]=8'h46;
    mem['h07D8]=8'h00; mem['h07D9]=8'h10; mem['h07DA]=8'h36; mem['h07DB]=8'h53;
    mem['h07DC]=8'h3E; mem['h07DD]=8'h00; mem['h07DE]=8'h44; mem['h07DF]=8'h34;
    mem['h07E0]=8'h10; mem['h07E1]=8'h36; mem['h07E2]=8'h0C; mem['h07E3]=8'h44;
    mem['h07E4]=8'hA4; mem['h07E5]=8'h12; mem['h07E6]=8'h36; mem['h07E7]=8'h56;
    mem['h07E8]=8'h2E; mem['h07E9]=8'h01; mem['h07EA]=8'hC7; mem['h07EB]=8'hA0;
    mem['h07EC]=8'h70; mem['h07ED]=8'h82; mem['h07EE]=8'h10; mem['h07EF]=8'h07;
    mem['h07F0]=8'h36; mem['h07F1]=8'h56; mem['h07F2]=8'h2E; mem['h07F3]=8'h01;
    mem['h07F4]=8'hC7; mem['h07F5]=8'hA0; mem['h07F6]=8'h2B; mem['h07F7]=8'h50;
    mem['h07F8]=8'hA2; mem['h07F9]=8'h06; mem['h07FA]=8'h36; mem['h07FB]=8'h14;
    mem['h07FC]=8'h44; mem['h07FD]=8'hA4; mem['h07FE]=8'h12; mem['h07FF]=8'h46;
    mem['h0800]=8'h00; mem['h0801]=8'h10; mem['h0802]=8'h36; mem['h0803]=8'h54;
    mem['h0804]=8'hC7; mem['h0805]=8'h46; mem['h0806]=8'h82; mem['h0807]=8'h03;
    mem['h0808]=8'h36; mem['h0809]=8'h7F; mem['h080A]=8'h2E; mem['h080B]=8'h16;
    mem['h080C]=8'h3E; mem['h080D]=8'hFF; mem['h080E]=8'h07; mem['h080F]=8'h46;
    mem['h0810]=8'h00; mem['h0811]=8'h10; mem['h0812]=8'h36; mem['h0813]=8'h54;
    mem['h0814]=8'hC7; mem['h0815]=8'h36; mem['h0816]=8'h23; mem['h0817]=8'h97;
    mem['h0818]=8'h36; mem['h0819]=8'h7F; mem['h081A]=8'h2E; mem['h081B]=8'h16;
    mem['h081C]=8'h3E; mem['h081D]=8'hFF; mem['h081E]=8'h70; mem['h081F]=8'h8F;
    mem['h0820]=8'h19; mem['h0821]=8'h2B; mem['h0822]=8'hD0; mem['h0823]=8'h06;
    mem['h0824]=8'hA0; mem['h0825]=8'h46; mem['h0826]=8'h82; mem['h0827]=8'h03;
    mem['h0828]=8'h11; mem['h0829]=8'h48; mem['h082A]=8'h25; mem['h082B]=8'h08;
    mem['h082C]=8'h07; mem['h082D]=8'h36; mem['h082E]=8'h81; mem['h082F]=8'h2E;
    mem['h0830]=8'h17; mem['h0831]=8'hC7; mem['h0832]=8'hA0; mem['h0833]=8'h68;
    mem['h0834]=8'h40; mem['h0835]=8'h08; mem['h0836]=8'h3E; mem['h0837]=8'h00;
    mem['h0838]=8'h36; mem['h0839]=8'h84; mem['h083A]=8'hF7; mem['h083B]=8'h2E;
    mem['h083C]=8'h2F; mem['h083D]=8'h44; mem['h083E]=8'hAD; mem['h083F]=8'h12;
    mem['h0840]=8'h36; mem['h0841]=8'hF8; mem['h0842]=8'h2E; mem['h0843]=8'h16;
    mem['h0844]=8'h3E; mem['h0845]=8'h00; mem['h0846]=8'h36; mem['h0847]=8'h50;
    mem['h0848]=8'h1E; mem['h0849]=8'h17; mem['h084A]=8'h26; mem['h084B]=8'h88;
    mem['h084C]=8'hC7; mem['h084D]=8'h3C; mem['h084E]=8'h01; mem['h084F]=8'h48;
    mem['h0850]=8'h56; mem['h0851]=8'h08; mem['h0852]=8'h36; mem['h0853]=8'h52;
    mem['h0854]=8'h3E; mem['h0855]=8'h00; mem['h0856]=8'h36; mem['h0857]=8'h51;
    mem['h0858]=8'h2E; mem['h0859]=8'h16; mem['h085A]=8'h46; mem['h085B]=8'hEE;
    mem['h085C]=8'h12; mem['h085D]=8'hC7; mem['h085E]=8'h30; mem['h085F]=8'hCF;
    mem['h0860]=8'h30; mem['h0861]=8'h46; mem['h0862]=8'hEE; mem['h0863]=8'h12;
    mem['h0864]=8'hBF; mem['h0865]=8'h48; mem['h0866]=8'h6E; mem['h0867]=8'h08;
    mem['h0868]=8'h30; mem['h0869]=8'hC1; mem['h086A]=8'hBF; mem['h086B]=8'h68;
    mem['h086C]=8'h97; mem['h086D]=8'h08; mem['h086E]=8'h46; mem['h086F]=8'hAE;
    mem['h0870]=8'h06; mem['h0871]=8'h36; mem['h0872]=8'hF8; mem['h0873]=8'h2E;
    mem['h0874]=8'h16; mem['h0875]=8'hCF; mem['h0876]=8'h08; mem['h0877]=8'hF9;
    mem['h0878]=8'h36; mem['h0879]=8'h3F; mem['h087A]=8'h2E; mem['h087B]=8'h17;
    mem['h087C]=8'hC1; mem['h087D]=8'hBF; mem['h087E]=8'h48; mem['h087F]=8'h56;
    mem['h0880]=8'h08; mem['h0881]=8'h36; mem['h0882]=8'h3F; mem['h0883]=8'h2E;
    mem['h0884]=8'h17; mem['h0885]=8'hCF; mem['h0886]=8'h08; mem['h0887]=8'hF9;
    mem['h0888]=8'hC1; mem['h0889]=8'h3C; mem['h088A]=8'h15; mem['h088B]=8'h50;
    mem['h088C]=8'h92; mem['h088D]=8'h02; mem['h088E]=8'h36; mem['h088F]=8'h51;
    mem['h0890]=8'h2E; mem['h0891]=8'h16; mem['h0892]=8'h0E; mem['h0893]=8'h02;
    mem['h0894]=8'h46; mem['h0895]=8'h0B; mem['h0896]=8'h11; mem['h0897]=8'h46;
    mem['h0898]=8'hEE; mem['h0899]=8'h12; mem['h089A]=8'h46; mem['h089B]=8'hAD;
    mem['h089C]=8'h12; mem['h089D]=8'h44; mem['h089E]=8'hAD; mem['h089F]=8'h02;
    mem['h08A0]=8'h36; mem['h08A1]=8'h50; mem['h08A2]=8'h2E; mem['h08A3]=8'h16;
    mem['h08A4]=8'hDD; mem['h08A5]=8'h26; mem['h08A6]=8'h64; mem['h08A7]=8'h44;
    mem['h08A8]=8'hB1; mem['h08A9]=8'h08; mem['h08AA]=8'h36; mem['h08AB]=8'h64;
    mem['h08AC]=8'h2E; mem['h08AD]=8'h16; mem['h08AE]=8'hDD; mem['h08AF]=8'h26;
    mem['h08B0]=8'h50; mem['h08B1]=8'hCF; mem['h08B2]=8'h08; mem['h08B3]=8'h44;
    mem['h08B4]=8'h0B; mem['h08B5]=8'h11; mem['h08B6]=8'h36; mem['h08B7]=8'hEA;
    mem['h08B8]=8'h2E; mem['h08B9]=8'h01; mem['h08BA]=8'h46; mem['h08BB]=8'h51;
    mem['h08BC]=8'h03; mem['h08BD]=8'h36; mem['h08BE]=8'h00; mem['h08BF]=8'h2E;
    mem['h08C0]=8'h16; mem['h08C1]=8'h46; mem['h08C2]=8'h0C; mem['h08C3]=8'h03;
    mem['h08C4]=8'hC7; mem['h08C5]=8'hA0; mem['h08C6]=8'h68; mem['h08C7]=8'hBD;
    mem['h08C8]=8'h08; mem['h08C9]=8'h36; mem['h08CA]=8'hDD; mem['h08CB]=8'h2E;
    mem['h08CC]=8'h01; mem['h08CD]=8'h1E; mem['h08CE]=8'h16; mem['h08CF]=8'h26;
    mem['h08D0]=8'h00; mem['h08D1]=8'h46; mem['h08D2]=8'hDA; mem['h08D3]=8'h02;
    mem['h08D4]=8'h48; mem['h08D5]=8'hEC; mem['h08D6]=8'h08; mem['h08D7]=8'h36;
    mem['h08D8]=8'h00; mem['h08D9]=8'h2E; mem['h08DA]=8'h1B; mem['h08DB]=8'hC7;
    mem['h08DC]=8'hA0; mem['h08DD]=8'h68; mem['h08DE]=8'hB6; mem['h08DF]=8'h08;
    mem['h08E0]=8'h46; mem['h08E1]=8'h51; mem['h08E2]=8'h03; mem['h08E3]=8'h46;
    mem['h08E4]=8'hFF; mem['h08E5]=8'h02; mem['h08E6]=8'h46; mem['h08E7]=8'h61;
    mem['h08E8]=8'h03; mem['h08E9]=8'h44; mem['h08EA]=8'hDB; mem['h08EB]=8'h08;
    mem['h08EC]=8'h36; mem['h08ED]=8'hE2; mem['h08EE]=8'h2E; mem['h08EF]=8'h01;
    mem['h08F0]=8'h26; mem['h08F1]=8'h00; mem['h08F2]=8'h1E; mem['h08F3]=8'h16;
    mem['h08F4]=8'h26; mem['h08F5]=8'h00; mem['h08F6]=8'h46; mem['h08F7]=8'hDA;
    mem['h08F8]=8'h02; mem['h08F9]=8'h68; mem['h08FA]=8'h38; mem['h08FB]=8'h0B;
    mem['h08FC]=8'h1E; mem['h08FD]=8'h16; mem['h08FE]=8'h26; mem['h08FF]=8'h00;
    mem['h0900]=8'h36; mem['h0901]=8'hE6; mem['h0902]=8'h2E; mem['h0903]=8'h01;
    mem['h0904]=8'h46; mem['h0905]=8'hDA; mem['h0906]=8'h02; mem['h0907]=8'h48;
    mem['h0908]=8'h39; mem['h0909]=8'h09; mem['h090A]=8'h2E; mem['h090B]=8'h16;
    mem['h090C]=8'h36; mem['h090D]=8'hF4; mem['h090E]=8'h3E; mem['h090F]=8'h1B;
    mem['h0910]=8'h30; mem['h0911]=8'h3E; mem['h0912]=8'h00; mem['h0913]=8'h36;
    mem['h0914]=8'h3F; mem['h0915]=8'h2E; mem['h0916]=8'h17; mem['h0917]=8'h3E;
    mem['h0918]=8'h01; mem['h0919]=8'h36; mem['h091A]=8'h3D; mem['h091B]=8'h3E;
    mem['h091C]=8'h00; mem['h091D]=8'h36; mem['h091E]=8'h50; mem['h091F]=8'h3E;
    mem['h0920]=8'h00; mem['h0921]=8'h36; mem['h0922]=8'h88; mem['h0923]=8'h3E;
    mem['h0924]=8'h00; mem['h0925]=8'h30; mem['h0926]=8'h3E; mem['h0927]=8'h00;
    mem['h0928]=8'h2E; mem['h0929]=8'h1B; mem['h092A]=8'h36; mem['h092B]=8'h00;
    mem['h092C]=8'h3E; mem['h092D]=8'h00; mem['h092E]=8'h2E; mem['h092F]=8'h2F;
    mem['h0930]=8'h3E; mem['h0931]=8'h00; mem['h0932]=8'h30; mem['h0933]=8'h48;
    mem['h0934]=8'h30; mem['h0935]=8'h09; mem['h0936]=8'h44; mem['h0937]=8'hB6;
    mem['h0938]=8'h08; mem['h0939]=8'h26; mem['h093A]=8'hBA; mem['h093B]=8'h1E;
    mem['h093C]=8'h01; mem['h093D]=8'h2E; mem['h093E]=8'h16; mem['h093F]=8'h36;
    mem['h0940]=8'h00; mem['h0941]=8'h46; mem['h0942]=8'hDA; mem['h0943]=8'h02;
    mem['h0944]=8'h68; mem['h0945]=8'h40; mem['h0946]=8'h00; mem['h0947]=8'h36;
    mem['h0948]=8'hBF; mem['h0949]=8'h2E; mem['h094A]=8'h01; mem['h094B]=8'h1E;
    mem['h094C]=8'h16; mem['h094D]=8'h26; mem['h094E]=8'h00; mem['h094F]=8'h46;
    mem['h0950]=8'hDA; mem['h0951]=8'h02; mem['h0952]=8'h68; mem['h0953]=8'h40;
    mem['h0954]=8'h00; mem['h0955]=8'h36; mem['h0956]=8'hF0; mem['h0957]=8'h2E;
    mem['h0958]=8'h16; mem['h0959]=8'h3E; mem['h095A]=8'h1B; mem['h095B]=8'h30;
    mem['h095C]=8'h3E; mem['h095D]=8'h00; mem['h095E]=8'h46; mem['h095F]=8'h00;
    mem['h0960]=8'h02; mem['h0961]=8'h36; mem['h0962]=8'h83; mem['h0963]=8'h2E;
    mem['h0964]=8'h16; mem['h0965]=8'hC7; mem['h0966]=8'hA0; mem['h0967]=8'h50;
    mem['h0968]=8'h71; mem['h0969]=8'h09; mem['h096A]=8'h06; mem['h096B]=8'hD3;
    mem['h096C]=8'h16; mem['h096D]=8'hD9; mem['h096E]=8'h44; mem['h096F]=8'h96;
    mem['h0970]=8'h02; mem['h0971]=8'h36; mem['h0972]=8'hE0; mem['h0973]=8'hC7;
    mem['h0974]=8'hA0; mem['h0975]=8'h68; mem['h0976]=8'h89; mem['h0977]=8'h0B;
    mem['h0978]=8'h36; mem['h0979]=8'hF0; mem['h097A]=8'h3E; mem['h097B]=8'h1B;
    mem['h097C]=8'h30; mem['h097D]=8'h3E; mem['h097E]=8'h00; mem['h097F]=8'h36;
    mem['h0980]=8'h81; mem['h0981]=8'h2E; mem['h0982]=8'h16; mem['h0983]=8'h3E;
    mem['h0984]=8'h01; mem['h0985]=8'h36; mem['h0986]=8'hE8; mem['h0987]=8'h3E;
    mem['h0988]=8'h00; mem['h0989]=8'h36; mem['h098A]=8'h81; mem['h098B]=8'h46;
    mem['h098C]=8'h53; mem['h098D]=8'h0A; mem['h098E]=8'h68; mem['h098F]=8'hA2;
    mem['h0990]=8'h09; mem['h0991]=8'h3C; mem['h0992]=8'hB0; mem['h0993]=8'h70;
    mem['h0994]=8'hB7; mem['h0995]=8'h09; mem['h0996]=8'h3C; mem['h0997]=8'hBA;
    mem['h0998]=8'h50; mem['h0999]=8'hB7; mem['h099A]=8'h09; mem['h099B]=8'h36;
    mem['h099C]=8'hE8; mem['h099D]=8'h2E; mem['h099E]=8'h16; mem['h099F]=8'h46;
    mem['h09A0]=8'hCC; mem['h09A1]=8'h02; mem['h09A2]=8'h36; mem['h09A3]=8'h81;
    mem['h09A4]=8'h2E; mem['h09A5]=8'h16; mem['h09A6]=8'hCF; mem['h09A7]=8'h08;
    mem['h09A8]=8'hF9; mem['h09A9]=8'h36; mem['h09AA]=8'hF0; mem['h09AB]=8'h2E;
    mem['h09AC]=8'h16; mem['h09AD]=8'hD7; mem['h09AE]=8'h30; mem['h09AF]=8'hF7;
    mem['h09B0]=8'hEA; mem['h09B1]=8'hC7; mem['h09B2]=8'h09; mem['h09B3]=8'hB9;
    mem['h09B4]=8'h48; mem['h09B5]=8'h89; mem['h09B6]=8'h09; mem['h09B7]=8'h36;
    mem['h09B8]=8'hF0; mem['h09B9]=8'h2E; mem['h09BA]=8'h16; mem['h09BB]=8'hDF;
    mem['h09BC]=8'h30; mem['h09BD]=8'hF7; mem['h09BE]=8'hEB; mem['h09BF]=8'hC7;
    mem['h09C0]=8'hA0; mem['h09C1]=8'h48; mem['h09C2]=8'hDE; mem['h09C3]=8'h09;
    mem['h09C4]=8'h44; mem['h09C5]=8'h05; mem['h09C6]=8'h0A; mem['h09C7]=8'h36;
    mem['h09C8]=8'h81; mem['h09C9]=8'h2E; mem['h09CA]=8'h17; mem['h09CB]=8'h3E;
    mem['h09CC]=8'h00; mem['h09CD]=8'h44; mem['h09CE]=8'hB6; mem['h09CF]=8'h08;
    mem['h09D0]=8'hFF; mem['h09D1]=8'hFF; mem['h09D2]=8'hFF; mem['h09D3]=8'hFF;
    mem['h09D4]=8'hFF; mem['h09D5]=8'hFF; mem['h09D6]=8'hFF; mem['h09D7]=8'hFF;
    mem['h09D8]=8'hFF; mem['h09D9]=8'hFF; mem['h09DA]=8'hFF; mem['h09DB]=8'hFF;
    mem['h09DC]=8'hFF; mem['h09DD]=8'hFF; mem['h09DE]=8'h36; mem['h09DF]=8'hE8;
    mem['h09E0]=8'h2E; mem['h09E1]=8'h16; mem['h09E2]=8'h1E; mem['h09E3]=8'h16;
    mem['h09E4]=8'h26; mem['h09E5]=8'hE0; mem['h09E6]=8'h46; mem['h09E7]=8'hDA;
    mem['h09E8]=8'h02; mem['h09E9]=8'h70; mem['h09EA]=8'h3B; mem['h09EB]=8'h0A;
    mem['h09EC]=8'h48; mem['h09ED]=8'h05; mem['h09EE]=8'h0A; mem['h09EF]=8'h36;
    mem['h09F0]=8'hF0; mem['h09F1]=8'h2E; mem['h09F2]=8'h16; mem['h09F3]=8'hD7;
    mem['h09F4]=8'h30; mem['h09F5]=8'hF7; mem['h09F6]=8'hEA; mem['h09F7]=8'hCF;
    mem['h09F8]=8'h08; mem['h09F9]=8'h46; mem['h09FA]=8'h64; mem['h09FB]=8'h0A;
    mem['h09FC]=8'h36; mem['h09FD]=8'h83; mem['h09FE]=8'h2E; mem['h09FF]=8'h16;
    mem['h0A00]=8'hC7; mem['h0A01]=8'hA0; mem['h0A02]=8'h68; mem['h0A03]=8'hB6;
    mem['h0A04]=8'h08; mem['h0A05]=8'h36; mem['h0A06]=8'hF0; mem['h0A07]=8'h2E;
    mem['h0A08]=8'h16; mem['h0A09]=8'hDF; mem['h0A0A]=8'h30; mem['h0A0B]=8'hE7;
    mem['h0A0C]=8'h36; mem['h0A0D]=8'h00; mem['h0A0E]=8'h2E; mem['h0A0F]=8'h16;
    mem['h0A10]=8'hCF; mem['h0A11]=8'h08; mem['h0A12]=8'h46; mem['h0A13]=8'h85;
    mem['h0A14]=8'h0A; mem['h0A15]=8'h36; mem['h0A16]=8'hF0; mem['h0A17]=8'h2E;
    mem['h0A18]=8'h16; mem['h0A19]=8'hDF; mem['h0A1A]=8'h30; mem['h0A1B]=8'hE7;
    mem['h0A1C]=8'h36; mem['h0A1D]=8'h00; mem['h0A1E]=8'h2E; mem['h0A1F]=8'h16;
    mem['h0A20]=8'h46; mem['h0A21]=8'h26; mem['h0A22]=8'h0A; mem['h0A23]=8'h44;
    mem['h0A24]=8'hBD; mem['h0A25]=8'h08; mem['h0A26]=8'hCF; mem['h0A27]=8'h08;
    mem['h0A28]=8'hC7; mem['h0A29]=8'h46; mem['h0A2A]=8'hFF; mem['h0A2B]=8'h02;
    mem['h0A2C]=8'h46; mem['h0A2D]=8'hEE; mem['h0A2E]=8'h12; mem['h0A2F]=8'hF8;
    mem['h0A30]=8'h46; mem['h0A31]=8'hFF; mem['h0A32]=8'h02; mem['h0A33]=8'h46;
    mem['h0A34]=8'hEE; mem['h0A35]=8'h12; mem['h0A36]=8'h09; mem['h0A37]=8'h48;
    mem['h0A38]=8'h28; mem['h0A39]=8'h0A; mem['h0A3A]=8'h07; mem['h0A3B]=8'h36;
    mem['h0A3C]=8'hF0; mem['h0A3D]=8'h2E; mem['h0A3E]=8'h16; mem['h0A3F]=8'hDF;
    mem['h0A40]=8'h30; mem['h0A41]=8'hE7; mem['h0A42]=8'hEB; mem['h0A43]=8'hF4;
    mem['h0A44]=8'hCF; mem['h0A45]=8'h08; mem['h0A46]=8'h46; mem['h0A47]=8'hC5;
    mem['h0A48]=8'h0A; mem['h0A49]=8'h36; mem['h0A4A]=8'hF0; mem['h0A4B]=8'h2E;
    mem['h0A4C]=8'h16; mem['h0A4D]=8'hFB; mem['h0A4E]=8'h30; mem['h0A4F]=8'hFC;
    mem['h0A50]=8'h44; mem['h0A51]=8'h7F; mem['h0A52]=8'h09; mem['h0A53]=8'h2E;
    mem['h0A54]=8'h16; mem['h0A55]=8'hCF; mem['h0A56]=8'h36; mem['h0A57]=8'hF0;
    mem['h0A58]=8'hDF; mem['h0A59]=8'h30; mem['h0A5A]=8'hE7; mem['h0A5B]=8'h46;
    mem['h0A5C]=8'hC5; mem['h0A5D]=8'h0A; mem['h0A5E]=8'hEB; mem['h0A5F]=8'hF4;
    mem['h0A60]=8'hC7; mem['h0A61]=8'h3C; mem['h0A62]=8'hA0; mem['h0A63]=8'h07;
    mem['h0A64]=8'h46; mem['h0A65]=8'h7C; mem['h0A66]=8'h03; mem['h0A67]=8'hD7;
    mem['h0A68]=8'h46; mem['h0A69]=8'h4B; mem['h0A6A]=8'h03; mem['h0A6B]=8'hFA;
    mem['h0A6C]=8'hC2; mem['h0A6D]=8'hA0; mem['h0A6E]=8'h68; mem['h0A6F]=8'h77;
    mem['h0A70]=8'h0A; mem['h0A71]=8'h46; mem['h0A72]=8'hFF; mem['h0A73]=8'h02;
    mem['h0A74]=8'h44; mem['h0A75]=8'h64; mem['h0A76]=8'h0A; mem['h0A77]=8'h36;
    mem['h0A78]=8'hF4; mem['h0A79]=8'h2E; mem['h0A7A]=8'h16; mem['h0A7B]=8'hDF;
    mem['h0A7C]=8'h30; mem['h0A7D]=8'hC7; mem['h0A7E]=8'h91; mem['h0A7F]=8'hF8;
    mem['h0A80]=8'h03; mem['h0A81]=8'h31; mem['h0A82]=8'h19; mem['h0A83]=8'hFB;
    mem['h0A84]=8'h07; mem['h0A85]=8'h36; mem['h0A86]=8'hF4; mem['h0A87]=8'h2E;
    mem['h0A88]=8'h16; mem['h0A89]=8'hC7; mem['h0A8A]=8'h30; mem['h0A8B]=8'hF7;
    mem['h0A8C]=8'hE8; mem['h0A8D]=8'h46; mem['h0A8E]=8'h7C; mem['h0A8F]=8'h03;
    mem['h0A90]=8'hC5; mem['h0A91]=8'h3C; mem['h0A92]=8'h2D; mem['h0A93]=8'h50;
    mem['h0A94]=8'h92; mem['h0A95]=8'h02; mem['h0A96]=8'h46; mem['h0A97]=8'h4B;
    mem['h0A98]=8'h03; mem['h0A99]=8'hD7; mem['h0A9A]=8'h46; mem['h0A9B]=8'h7C;
    mem['h0A9C]=8'h03; mem['h0A9D]=8'hFA; mem['h0A9E]=8'h46; mem['h0A9F]=8'h4B;
    mem['h0AA0]=8'h03; mem['h0AA1]=8'h46; mem['h0AA2]=8'hBF; mem['h0AA3]=8'h0A;
    mem['h0AA4]=8'h68; mem['h0AA5]=8'hAD; mem['h0AA6]=8'h0A; mem['h0AA7]=8'h46;
    mem['h0AA8]=8'h74; mem['h0AA9]=8'h03; mem['h0AAA]=8'h44; mem['h0AAB]=8'h99;
    mem['h0AAC]=8'h0A; mem['h0AAD]=8'h36; mem['h0AAE]=8'h00; mem['h0AAF]=8'h2E;
    mem['h0AB0]=8'h16; mem['h0AB1]=8'hCF; mem['h0AB2]=8'h08; mem['h0AB3]=8'h36;
    mem['h0AB4]=8'hF4; mem['h0AB5]=8'hDF; mem['h0AB6]=8'h30; mem['h0AB7]=8'hE7;
    mem['h0AB8]=8'h46; mem['h0AB9]=8'hC5; mem['h0ABA]=8'h0A; mem['h0ABB]=8'hFC;
    mem['h0ABC]=8'h31; mem['h0ABD]=8'hFB; mem['h0ABE]=8'h07; mem['h0ABF]=8'hC5;
    mem['h0AC0]=8'hBB; mem['h0AC1]=8'h0B; mem['h0AC2]=8'hC6; mem['h0AC3]=8'hBC;
    mem['h0AC4]=8'h07; mem['h0AC5]=8'hC4; mem['h0AC6]=8'h81; mem['h0AC7]=8'hE0;
    mem['h0AC8]=8'h03; mem['h0AC9]=8'h18; mem['h0ACA]=8'h07; mem['h0ACB]=8'h06;
    mem['h0ACC]=8'hDE; mem['h0ACD]=8'h16; mem['h0ACE]=8'hC3; mem['h0ACF]=8'h44;
    mem['h0AD0]=8'h96; mem['h0AD1]=8'h02; mem['h0AD2]=8'h36; mem['h0AD3]=8'hE0;
    mem['h0AD4]=8'h2E; mem['h0AD5]=8'h16; mem['h0AD6]=8'hC7; mem['h0AD7]=8'hA0;
    mem['h0AD8]=8'h68; mem['h0AD9]=8'hE9; mem['h0ADA]=8'h0A; mem['h0ADB]=8'h36;
    mem['h0ADC]=8'hF6; mem['h0ADD]=8'h2E; mem['h0ADE]=8'h01; mem['h0ADF]=8'h46;
    mem['h0AE0]=8'h51; mem['h0AE1]=8'h03; mem['h0AE2]=8'h36; mem['h0AE3]=8'hE0;
    mem['h0AE4]=8'h2E; mem['h0AE5]=8'h16; mem['h0AE6]=8'h46; mem['h0AE7]=8'h51;
    mem['h0AE8]=8'h03; mem['h0AE9]=8'h46; mem['h0AEA]=8'h61; mem['h0AEB]=8'h03;
    mem['h0AEC]=8'h44; mem['h0AED]=8'hC7; mem['h0AEE]=8'h09; mem['h0AEF]=8'h06;
    mem['h0AF0]=8'hC4; mem['h0AF1]=8'h16; mem['h0AF2]=8'hDA; mem['h0AF3]=8'h44;
    mem['h0AF4]=8'h96; mem['h0AF5]=8'h02; mem['h0AF6]=8'h06; mem['h0AF7]=8'hC6;
    mem['h0AF8]=8'h16; mem['h0AF9]=8'hD8; mem['h0AFA]=8'h44; mem['h0AFB]=8'h96;
    mem['h0AFC]=8'h02; mem['h0AFD]=8'h06; mem['h0AFE]=8'hC9; mem['h0AFF]=8'h16;
    mem['h0B00]=8'hCE; mem['h0B01]=8'h36; mem['h0B02]=8'h90; mem['h0B03]=8'h2E;
    mem['h0B04]=8'h01; mem['h0B05]=8'h3E; mem['h0B06]=8'h00; mem['h0B07]=8'h44;
    mem['h0B08]=8'h96; mem['h0B09]=8'h02; mem['h0B0A]=8'h1E; mem['h0B0B]=8'h16;
    mem['h0B0C]=8'h26; mem['h0B0D]=8'h00; mem['h0B0E]=8'h46; mem['h0B0F]=8'h34;
    mem['h0B10]=8'h0B; mem['h0B11]=8'h46; mem['h0B12]=8'hCF; mem['h0B13]=8'h12;
    mem['h0B14]=8'hCF; mem['h0B15]=8'h46; mem['h0B16]=8'hFF; mem['h0B17]=8'h02;
    mem['h0B18]=8'h46; mem['h0B19]=8'hF8; mem['h0B1A]=8'h02; mem['h0B1B]=8'h68;
    mem['h0B1C]=8'hDF; mem['h0B1D]=8'h12; mem['h0B1E]=8'h46; mem['h0B1F]=8'hDF;
    mem['h0B20]=8'h12; mem['h0B21]=8'h36; mem['h0B22]=8'h00; mem['h0B23]=8'h2E;
    mem['h0B24]=8'h16; mem['h0B25]=8'hC7; mem['h0B26]=8'hBC; mem['h0B27]=8'h68;
    mem['h0B28]=8'h31; mem['h0B29]=8'h0B; mem['h0B2A]=8'h46; mem['h0B2B]=8'hDF;
    mem['h0B2C]=8'h12; mem['h0B2D]=8'h44; mem['h0B2E]=8'h0E; mem['h0B2F]=8'h0B;
    mem['h0B30]=8'h00; mem['h0B31]=8'h26; mem['h0B32]=8'h00; mem['h0B33]=8'h07;
    mem['h0B34]=8'h20; mem['h0B35]=8'h0B; mem['h0B36]=8'h18; mem['h0B37]=8'h07;
    mem['h0B38]=8'h36; mem['h0B39]=8'h3B; mem['h0B3A]=8'h2E; mem['h0B3B]=8'h17;
    mem['h0B3C]=8'h3E; mem['h0B3D]=8'h00; mem['h0B3E]=8'h36; mem['h0B3F]=8'h85;
    mem['h0B40]=8'h3E; mem['h0B41]=8'h00; mem['h0B42]=8'h36; mem['h0B43]=8'hF0;
    mem['h0B44]=8'h2E; mem['h0B45]=8'h16; mem['h0B46]=8'h3E; mem['h0B47]=8'h1B;
    mem['h0B48]=8'h30; mem['h0B49]=8'h3E; mem['h0B4A]=8'h00; mem['h0B4B]=8'h44;
    mem['h0B4C]=8'h6E; mem['h0B4D]=8'h0B; mem['h0B4E]=8'h36; mem['h0B4F]=8'hF0;
    mem['h0B50]=8'h2E; mem['h0B51]=8'h16; mem['h0B52]=8'hDF; mem['h0B53]=8'h30;
    mem['h0B54]=8'hE7; mem['h0B55]=8'hEB; mem['h0B56]=8'hF4; mem['h0B57]=8'hCF;
    mem['h0B58]=8'h08; mem['h0B59]=8'h46; mem['h0B5A]=8'hC5; mem['h0B5B]=8'h0A;
    mem['h0B5C]=8'h36; mem['h0B5D]=8'hF0; mem['h0B5E]=8'h2E; mem['h0B5F]=8'h16;
    mem['h0B60]=8'hFB; mem['h0B61]=8'h30; mem['h0B62]=8'hFC; mem['h0B63]=8'h36;
    mem['h0B64]=8'hE0; mem['h0B65]=8'h2E; mem['h0B66]=8'h16; mem['h0B67]=8'hC7;
    mem['h0B68]=8'hA0; mem['h0B69]=8'h68; mem['h0B6A]=8'hB6; mem['h0B6B]=8'h08;
    mem['h0B6C]=8'hC0; mem['h0B6D]=8'hC0; mem['h0B6E]=8'h36; mem['h0B6F]=8'hF0;
    mem['h0B70]=8'h2E; mem['h0B71]=8'h16; mem['h0B72]=8'hD7; mem['h0B73]=8'h30;
    mem['h0B74]=8'hF7; mem['h0B75]=8'hEA; mem['h0B76]=8'h1E; mem['h0B77]=8'h16;
    mem['h0B78]=8'h26; mem['h0B79]=8'h00; mem['h0B7A]=8'h46; mem['h0B7B]=8'h26;
    mem['h0B7C]=8'h0A; mem['h0B7D]=8'h36; mem['h0B7E]=8'h00; mem['h0B7F]=8'h2E;
    mem['h0B80]=8'h16; mem['h0B81]=8'hC7; mem['h0B82]=8'hA0; mem['h0B83]=8'h68;
    mem['h0B84]=8'hB6; mem['h0B85]=8'h08; mem['h0B86]=8'h46; mem['h0B87]=8'h00;
    mem['h0B88]=8'h02; mem['h0B89]=8'h36; mem['h0B8A]=8'h83; mem['h0B8B]=8'h2E;
    mem['h0B8C]=8'h16; mem['h0B8D]=8'hC7; mem['h0B8E]=8'h3C; mem['h0B8F]=8'h01;
    mem['h0B90]=8'h68; mem['h0B91]=8'h4E; mem['h0B92]=8'h0B; mem['h0B93]=8'h3C;
    mem['h0B94]=8'h02; mem['h0B95]=8'h68; mem['h0B96]=8'h17; mem['h0B97]=8'h0E;
    mem['h0B98]=8'h3C; mem['h0B99]=8'h03; mem['h0B9A]=8'h68; mem['h0B9B]=8'h19;
    mem['h0B9C]=8'h0D; mem['h0B9D]=8'h3C; mem['h0B9E]=8'h04; mem['h0B9F]=8'h68;
    mem['h0BA0]=8'h7C; mem['h0BA1]=8'h0D; mem['h0BA2]=8'h3C; mem['h0BA3]=8'h05;
    mem['h0BA4]=8'h68; mem['h0BA5]=8'hE5; mem['h0BA6]=8'h0B; mem['h0BA7]=8'h3C;
    mem['h0BA8]=8'h06; mem['h0BA9]=8'h68; mem['h0BAA]=8'hF5; mem['h0BAB]=8'h0E;
    mem['h0BAC]=8'h3C; mem['h0BAD]=8'h07; mem['h0BAE]=8'h68; mem['h0BAF]=8'h74;
    mem['h0BB0]=8'h0F; mem['h0BB1]=8'h3C; mem['h0BB2]=8'h08; mem['h0BB3]=8'h68;
    mem['h0BB4]=8'h0B; mem['h0BB5]=8'h18; mem['h0BB6]=8'h3C; mem['h0BB7]=8'h09;
    mem['h0BB8]=8'h68; mem['h0BB9]=8'h9E; mem['h0BBA]=8'h0E; mem['h0BBB]=8'h3C;
    mem['h0BBC]=8'h0A; mem['h0BBD]=8'h68; mem['h0BBE]=8'hC4; mem['h0BBF]=8'h0E;
    mem['h0BC0]=8'h3C; mem['h0BC1]=8'h0B; mem['h0BC2]=8'h68; mem['h0BC3]=8'hF5;
    mem['h0BC4]=8'h2D; mem['h0BC5]=8'h3C; mem['h0BC6]=8'h0C; mem['h0BC7]=8'h68;
    mem['h0BC8]=8'hB6; mem['h0BC9]=8'h08; mem['h0BCA]=8'h3C; mem['h0BCB]=8'h0D;
    mem['h0BCC]=8'h68; mem['h0BCD]=8'h0B; mem['h0BCE]=8'h0D; mem['h0BCF]=8'h3C;
    mem['h0BD0]=8'h0E; mem['h0BD1]=8'h48; mem['h0BD2]=8'h6A; mem['h0BD3]=8'h09;
    mem['h0BD4]=8'h46; mem['h0BD5]=8'h6B; mem['h0BD6]=8'h2D; mem['h0BD7]=8'h36;
    mem['h0BD8]=8'h86; mem['h0BD9]=8'h2E; mem['h0BDA]=8'h16; mem['h0BDB]=8'hCF;
    mem['h0BDC]=8'h36; mem['h0BDD]=8'h82; mem['h0BDE]=8'hF9; mem['h0BDF]=8'h46;
    mem['h0BE0]=8'hA0; mem['h0BE1]=8'h08; mem['h0BE2]=8'h44; mem['h0BE3]=8'h22;
    mem['h0BE4]=8'h0D; mem['h0BE5]=8'h36; mem['h0BE6]=8'h82; mem['h0BE7]=8'h2E;
    mem['h0BE8]=8'h16; mem['h0BE9]=8'hC7; mem['h0BEA]=8'h36; mem['h0BEB]=8'h00;
    mem['h0BEC]=8'hBF; mem['h0BED]=8'h70; mem['h0BEE]=8'hF6; mem['h0BEF]=8'h0B;
    mem['h0BF0]=8'h46; mem['h0BF1]=8'h61; mem['h0BF2]=8'h03; mem['h0BF3]=8'h44;
    mem['h0BF4]=8'h4E; mem['h0BF5]=8'h0B; mem['h0BF6]=8'h46; mem['h0BF7]=8'hAD;
    mem['h0BF8]=8'h02; mem['h0BF9]=8'h36; mem['h0BFA]=8'h82; mem['h0BFB]=8'h2E;
    mem['h0BFC]=8'h16; mem['h0BFD]=8'hCF; mem['h0BFE]=8'h08; mem['h0BFF]=8'h36;
    mem['h0C00]=8'h83; mem['h0C01]=8'hF9; mem['h0C02]=8'h36; mem['h0C03]=8'h83;
    mem['h0C04]=8'h46; mem['h0C05]=8'hA0; mem['h0C06]=8'h02; mem['h0C07]=8'h3C;
    mem['h0C08]=8'hA7; mem['h0C09]=8'h68; mem['h0C0A]=8'h83; mem['h0C0B]=8'h0C;
    mem['h0C0C]=8'h3C; mem['h0C0D]=8'hA2; mem['h0C0E]=8'h68; mem['h0C0F]=8'h83;
    mem['h0C10]=8'h0C; mem['h0C11]=8'h3C; mem['h0C12]=8'hAC; mem['h0C13]=8'h68;
    mem['h0C14]=8'h23; mem['h0C15]=8'h0C; mem['h0C16]=8'h3C; mem['h0C17]=8'hBB;
    mem['h0C18]=8'h68; mem['h0C19]=8'h23; mem['h0C1A]=8'h0C; mem['h0C1B]=8'h36;
    mem['h0C1C]=8'h83; mem['h0C1D]=8'h46; mem['h0C1E]=8'h03; mem['h0C1F]=8'h03;
    mem['h0C20]=8'h48; mem['h0C21]=8'h02; mem['h0C22]=8'h0C; mem['h0C23]=8'h36;
    mem['h0C24]=8'h82; mem['h0C25]=8'hCF; mem['h0C26]=8'h08; mem['h0C27]=8'h36;
    mem['h0C28]=8'hBE; mem['h0C29]=8'hF9; mem['h0C2A]=8'h36; mem['h0C2B]=8'h83;
    mem['h0C2C]=8'hCF; mem['h0C2D]=8'h09; mem['h0C2E]=8'h36; mem['h0C2F]=8'hBF;
    mem['h0C30]=8'hF9; mem['h0C31]=8'h36; mem['h0C32]=8'hF7; mem['h0C33]=8'hC7;
    mem['h0C34]=8'hA0; mem['h0C35]=8'h68; mem['h0C36]=8'h3D; mem['h0C37]=8'h0C;
    mem['h0C38]=8'h3E; mem['h0C39]=8'h00; mem['h0C3A]=8'h44; mem['h0C3B]=8'h55;
    mem['h0C3C]=8'h0C; mem['h0C3D]=8'h46; mem['h0C3E]=8'h94; mem['h0C3F]=8'h03;
    mem['h0C40]=8'h36; mem['h0C41]=8'h7F; mem['h0C42]=8'h2E; mem['h0C43]=8'h16;
    mem['h0C44]=8'hC7; mem['h0C45]=8'hA0; mem['h0C46]=8'h36; mem['h0C47]=8'h48;
    mem['h0C48]=8'h2E; mem['h0C49]=8'h01; mem['h0C4A]=8'h3E; mem['h0C4B]=8'hFF;
    mem['h0C4C]=8'h6A; mem['h0C4D]=8'hCC; mem['h0C4E]=8'h0C; mem['h0C4F]=8'h36;
    mem['h0C50]=8'h7F; mem['h0C51]=8'h2E; mem['h0C52]=8'h16; mem['h0C53]=8'h3E;
    mem['h0C54]=8'h00; mem['h0C55]=8'h36; mem['h0C56]=8'h83; mem['h0C57]=8'h46;
    mem['h0C58]=8'hA0; mem['h0C59]=8'h02; mem['h0C5A]=8'h3C; mem['h0C5B]=8'hAC;
    mem['h0C5C]=8'h6A; mem['h0C5D]=8'hEF; mem['h0C5E]=8'h0C; mem['h0C5F]=8'h36;
    mem['h0C60]=8'h83; mem['h0C61]=8'h2E; mem['h0C62]=8'h16; mem['h0C63]=8'hCF;
    mem['h0C64]=8'h36; mem['h0C65]=8'h82; mem['h0C66]=8'hF9; mem['h0C67]=8'h36;
    mem['h0C68]=8'h00; mem['h0C69]=8'hC1; mem['h0C6A]=8'hBF; mem['h0C6B]=8'h70;
    mem['h0C6C]=8'hF6; mem['h0C6D]=8'h0B; mem['h0C6E]=8'h36; mem['h0C6F]=8'h00;
    mem['h0C70]=8'h46; mem['h0C71]=8'hA0; mem['h0C72]=8'h02; mem['h0C73]=8'h3C;
    mem['h0C74]=8'hAC; mem['h0C75]=8'h68; mem['h0C76]=8'h4E; mem['h0C77]=8'h0B;
    mem['h0C78]=8'h3C; mem['h0C79]=8'hBB; mem['h0C7A]=8'h68; mem['h0C7B]=8'h4E;
    mem['h0C7C]=8'h0B; mem['h0C7D]=8'h46; mem['h0C7E]=8'h61; mem['h0C7F]=8'h03;
    mem['h0C80]=8'h44; mem['h0C81]=8'h4E; mem['h0C82]=8'h0B; mem['h0C83]=8'h36;
    mem['h0C84]=8'hF7; mem['h0C85]=8'hF8; mem['h0C86]=8'h46; mem['h0C87]=8'hAD;
    mem['h0C88]=8'h02; mem['h0C89]=8'h36; mem['h0C8A]=8'h83; mem['h0C8B]=8'hCF;
    mem['h0C8C]=8'h08; mem['h0C8D]=8'h36; mem['h0C8E]=8'h84; mem['h0C8F]=8'hF9;
    mem['h0C90]=8'h36; mem['h0C91]=8'h84; mem['h0C92]=8'h46; mem['h0C93]=8'hA0;
    mem['h0C94]=8'h02; mem['h0C95]=8'h36; mem['h0C96]=8'hF7; mem['h0C97]=8'hBF;
    mem['h0C98]=8'h68; mem['h0C99]=8'hB3; mem['h0C9A]=8'h0C; mem['h0C9B]=8'h46;
    mem['h0C9C]=8'h82; mem['h0C9D]=8'h03; mem['h0C9E]=8'h36; mem['h0C9F]=8'h84;
    mem['h0CA0]=8'h46; mem['h0CA1]=8'h03; mem['h0CA2]=8'h03; mem['h0CA3]=8'h48;
    mem['h0CA4]=8'h90; mem['h0CA5]=8'h0C; mem['h0CA6]=8'h06; mem['h0CA7]=8'hC9;
    mem['h0CA8]=8'h16; mem['h0CA9]=8'hD1; mem['h0CAA]=8'h36; mem['h0CAB]=8'hF7;
    mem['h0CAC]=8'h2E; mem['h0CAD]=8'h16; mem['h0CAE]=8'h3E; mem['h0CAF]=8'h00;
    mem['h0CB0]=8'h44; mem['h0CB1]=8'h96; mem['h0CB2]=8'h02; mem['h0CB3]=8'h36;
    mem['h0CB4]=8'h84; mem['h0CB5]=8'hCF; mem['h0CB6]=8'h36; mem['h0CB7]=8'h82;
    mem['h0CB8]=8'hF9; mem['h0CB9]=8'hC1; mem['h0CBA]=8'h36; mem['h0CBB]=8'h00;
    mem['h0CBC]=8'hBF; mem['h0CBD]=8'h48; mem['h0CBE]=8'hF6; mem['h0CBF]=8'h0B;
    mem['h0CC0]=8'h46; mem['h0CC1]=8'h61; mem['h0CC2]=8'h03; mem['h0CC3]=8'h36;
    mem['h0CC4]=8'hF7; mem['h0CC5]=8'h2E; mem['h0CC6]=8'h16; mem['h0CC7]=8'h3E;
    mem['h0CC8]=8'h00; mem['h0CC9]=8'h44; mem['h0CCA]=8'h4E; mem['h0CCB]=8'h0B;
    mem['h0CCC]=8'h36; mem['h0CCD]=8'h56; mem['h0CCE]=8'h2E; mem['h0CCF]=8'h01;
    mem['h0CD0]=8'hC7; mem['h0CD1]=8'hA0; mem['h0CD2]=8'h68; mem['h0CD3]=8'hDE;
    mem['h0CD4]=8'h0C; mem['h0CD5]=8'h30; mem['h0CD6]=8'hC7; mem['h0CD7]=8'hA0;
    mem['h0CD8]=8'h68; mem['h0CD9]=8'hE8; mem['h0CDA]=8'h0C; mem['h0CDB]=8'h44;
    mem['h0CDC]=8'h75; mem['h0CDD]=8'h14; mem['h0CDE]=8'h06; mem['h0CDF]=8'hA0;
    mem['h0CE0]=8'h46; mem['h0CE1]=8'h82; mem['h0CE2]=8'h03; mem['h0CE3]=8'h06;
    mem['h0CE4]=8'hB0; mem['h0CE5]=8'h44; mem['h0CE6]=8'h82; mem['h0CE7]=8'h03;
    mem['h0CE8]=8'h36; mem['h0CE9]=8'h48; mem['h0CEA]=8'h3E; mem['h0CEB]=8'h00;
    mem['h0CEC]=8'h44; mem['h0CED]=8'h75; mem['h0CEE]=8'h14; mem['h0CEF]=8'h36;
    mem['h0CF0]=8'h00; mem['h0CF1]=8'hC7; mem['h0CF2]=8'h36; mem['h0CF3]=8'h83;
    mem['h0CF4]=8'h97; mem['h0CF5]=8'h33; mem['h0CF6]=8'h36; mem['h0CF7]=8'h23;
    mem['h0CF8]=8'h2E; mem['h0CF9]=8'h01; mem['h0CFA]=8'hC7; mem['h0CFB]=8'h24;
    mem['h0CFC]=8'hF0; mem['h0CFD]=8'h04; mem['h0CFE]=8'h10; mem['h0CFF]=8'h97;
    mem['h0D00]=8'hD0; mem['h0D01]=8'h06; mem['h0D02]=8'hA0; mem['h0D03]=8'h46;
    mem['h0D04]=8'h82; mem['h0D05]=8'h03; mem['h0D06]=8'h11; mem['h0D07]=8'h48;
    mem['h0D08]=8'h03; mem['h0D09]=8'h0D; mem['h0D0A]=8'h07; mem['h0D0B]=8'h46;
    mem['h0D0C]=8'hA0; mem['h0D0D]=8'h08; mem['h0D0E]=8'h36; mem['h0D0F]=8'h82;
    mem['h0D10]=8'h2E; mem['h0D11]=8'h16; mem['h0D12]=8'hCF; mem['h0D13]=8'h36;
    mem['h0D14]=8'h83; mem['h0D15]=8'hF9; mem['h0D16]=8'h44; mem['h0D17]=8'h61;
    mem['h0D18]=8'h0D; mem['h0D19]=8'h46; mem['h0D1A]=8'hAD; mem['h0D1B]=8'h02;
    mem['h0D1C]=8'h36; mem['h0D1D]=8'h64; mem['h0D1E]=8'h2E; mem['h0D1F]=8'h16;
    mem['h0D20]=8'h3E; mem['h0D21]=8'h00; mem['h0D22]=8'h36; mem['h0D23]=8'h82;
    mem['h0D24]=8'h2E; mem['h0D25]=8'h16; mem['h0D26]=8'hCF; mem['h0D27]=8'h08;
    mem['h0D28]=8'h36; mem['h0D29]=8'h83; mem['h0D2A]=8'hF9; mem['h0D2B]=8'h36;
    mem['h0D2C]=8'h83; mem['h0D2D]=8'h46; mem['h0D2E]=8'hA0; mem['h0D2F]=8'h02;
    mem['h0D30]=8'h68; mem['h0D31]=8'h52; mem['h0D32]=8'h0D; mem['h0D33]=8'h3C;
    mem['h0D34]=8'hBD; mem['h0D35]=8'h68; mem['h0D36]=8'h61; mem['h0D37]=8'h0D;
    mem['h0D38]=8'h3C; mem['h0D39]=8'hA8; mem['h0D3A]=8'h48; mem['h0D3B]=8'h4B;
    mem['h0D3C]=8'h0D; mem['h0D3D]=8'h46; mem['h0D3E]=8'h65; mem['h0D3F]=8'h2D;
    mem['h0D40]=8'h36; mem['h0D41]=8'h86; mem['h0D42]=8'h2E; mem['h0D43]=8'h16;
    mem['h0D44]=8'hCF; mem['h0D45]=8'h36; mem['h0D46]=8'h83; mem['h0D47]=8'hF9;
    mem['h0D48]=8'h44; mem['h0D49]=8'h52; mem['h0D4A]=8'h0D; mem['h0D4B]=8'h36;
    mem['h0D4C]=8'h64; mem['h0D4D]=8'h2E; mem['h0D4E]=8'h16; mem['h0D4F]=8'h46;
    mem['h0D50]=8'hCC; mem['h0D51]=8'h02; mem['h0D52]=8'h36; mem['h0D53]=8'h83;
    mem['h0D54]=8'h46; mem['h0D55]=8'h03; mem['h0D56]=8'h03; mem['h0D57]=8'h48;
    mem['h0D58]=8'h2B; mem['h0D59]=8'h0D; mem['h0D5A]=8'h06; mem['h0D5B]=8'hCC;
    mem['h0D5C]=8'h16; mem['h0D5D]=8'hC5; mem['h0D5E]=8'h44; mem['h0D5F]=8'h96;
    mem['h0D60]=8'h02; mem['h0D61]=8'h36; mem['h0D62]=8'h83; mem['h0D63]=8'h2E;
    mem['h0D64]=8'h16; mem['h0D65]=8'hCF; mem['h0D66]=8'h08; mem['h0D67]=8'h36;
    mem['h0D68]=8'hBE; mem['h0D69]=8'hF9; mem['h0D6A]=8'h36; mem['h0D6B]=8'h00;
    mem['h0D6C]=8'hCF; mem['h0D6D]=8'h36; mem['h0D6E]=8'hBF; mem['h0D6F]=8'hF9;
    mem['h0D70]=8'h46; mem['h0D71]=8'h94; mem['h0D72]=8'h03; mem['h0D73]=8'h46;
    mem['h0D74]=8'hAA; mem['h0D75]=8'h08; mem['h0D76]=8'h46; mem['h0D77]=8'h2D;
    mem['h0D78]=8'h08; mem['h0D79]=8'h44; mem['h0D7A]=8'h4E; mem['h0D7B]=8'h0B;
    mem['h0D7C]=8'h36; mem['h0D7D]=8'hE8; mem['h0D7E]=8'h2E; mem['h0D7F]=8'h16;
    mem['h0D80]=8'h3E; mem['h0D81]=8'h00; mem['h0D82]=8'h36; mem['h0D83]=8'h82;
    mem['h0D84]=8'hCF; mem['h0D85]=8'h08; mem['h0D86]=8'h36; mem['h0D87]=8'h83;
    mem['h0D88]=8'hF9; mem['h0D89]=8'h36; mem['h0D8A]=8'h83; mem['h0D8B]=8'h46;
    mem['h0D8C]=8'hA0; mem['h0D8D]=8'h02; mem['h0D8E]=8'h68; mem['h0D8F]=8'hA0;
    mem['h0D90]=8'h0D; mem['h0D91]=8'h3C; mem['h0D92]=8'hB0; mem['h0D93]=8'h70;
    mem['h0D94]=8'hA8; mem['h0D95]=8'h0D; mem['h0D96]=8'h3C; mem['h0D97]=8'hBA;
    mem['h0D98]=8'h50; mem['h0D99]=8'hA8; mem['h0D9A]=8'h0D; mem['h0D9B]=8'h36;
    mem['h0D9C]=8'hE8; mem['h0D9D]=8'h46; mem['h0D9E]=8'hCC; mem['h0D9F]=8'h02;
    mem['h0DA0]=8'h36; mem['h0DA1]=8'h83; mem['h0DA2]=8'h46; mem['h0DA3]=8'h03;
    mem['h0DA4]=8'h03; mem['h0DA5]=8'h48; mem['h0DA6]=8'h89; mem['h0DA7]=8'h0D;
    mem['h0DA8]=8'h36; mem['h0DA9]=8'hF0; mem['h0DAA]=8'h2E; mem['h0DAB]=8'h16;
    mem['h0DAC]=8'h3E; mem['h0DAD]=8'h1B; mem['h0DAE]=8'h30; mem['h0DAF]=8'h3E;
    mem['h0DB0]=8'h00; mem['h0DB1]=8'h46; mem['h0DB2]=8'hAD; mem['h0DB3]=8'h02;
    mem['h0DB4]=8'h36; mem['h0DB5]=8'h84; mem['h0DB6]=8'h3E; mem['h0DB7]=8'h01;
    mem['h0DB8]=8'h36; mem['h0DB9]=8'h84; mem['h0DBA]=8'h46; mem['h0DBB]=8'h53;
    mem['h0DBC]=8'h0A; mem['h0DBD]=8'h68; mem['h0DBE]=8'hCD; mem['h0DBF]=8'h0D;
    mem['h0DC0]=8'h3C; mem['h0DC1]=8'hB0; mem['h0DC2]=8'h70; mem['h0DC3]=8'hE0;
    mem['h0DC4]=8'h0D; mem['h0DC5]=8'h3C; mem['h0DC6]=8'hBA; mem['h0DC7]=8'h50;
    mem['h0DC8]=8'hE0; mem['h0DC9]=8'h0D; mem['h0DCA]=8'h46; mem['h0DCB]=8'hC8;
    mem['h0DCC]=8'h02; mem['h0DCD]=8'h36; mem['h0DCE]=8'h84; mem['h0DCF]=8'h2E;
    mem['h0DD0]=8'h16; mem['h0DD1]=8'hCF; mem['h0DD2]=8'h08; mem['h0DD3]=8'hF9;
    mem['h0DD4]=8'h36; mem['h0DD5]=8'hF0; mem['h0DD6]=8'hD7; mem['h0DD7]=8'h30;
    mem['h0DD8]=8'hF7; mem['h0DD9]=8'hEA; mem['h0DDA]=8'hC7; mem['h0DDB]=8'h09;
    mem['h0DDC]=8'hB9; mem['h0DDD]=8'h48; mem['h0DDE]=8'hB8; mem['h0DDF]=8'h0D;
    mem['h0DE0]=8'h36; mem['h0DE1]=8'h50; mem['h0DE2]=8'h2E; mem['h0DE3]=8'h16;
    mem['h0DE4]=8'h1E; mem['h0DE5]=8'h16; mem['h0DE6]=8'h26; mem['h0DE7]=8'hE8;
    mem['h0DE8]=8'h46; mem['h0DE9]=8'hDA; mem['h0DEA]=8'h02; mem['h0DEB]=8'h68;
    mem['h0DEC]=8'h6E; mem['h0DED]=8'h0B; mem['h0DEE]=8'h36; mem['h0DEF]=8'hF0;
    mem['h0DF0]=8'h2E; mem['h0DF1]=8'h16; mem['h0DF2]=8'hDF; mem['h0DF3]=8'h30;
    mem['h0DF4]=8'hE7; mem['h0DF5]=8'hEB; mem['h0DF6]=8'hF4; mem['h0DF7]=8'hCF;
    mem['h0DF8]=8'h08; mem['h0DF9]=8'h46; mem['h0DFA]=8'hC5; mem['h0DFB]=8'h0A;
    mem['h0DFC]=8'h36; mem['h0DFD]=8'hF0; mem['h0DFE]=8'h2E; mem['h0DFF]=8'h16;
    mem['h0E00]=8'hFB; mem['h0E01]=8'h30; mem['h0E02]=8'hFC; mem['h0E03]=8'h36;
    mem['h0E04]=8'hF4; mem['h0E05]=8'hC3; mem['h0E06]=8'hBF; mem['h0E07]=8'h48;
    mem['h0E08]=8'hB1; mem['h0E09]=8'h0D; mem['h0E0A]=8'h30; mem['h0E0B]=8'hC4;
    mem['h0E0C]=8'hBF; mem['h0E0D]=8'h48; mem['h0E0E]=8'hB1; mem['h0E0F]=8'h0D;
    mem['h0E10]=8'h06; mem['h0E11]=8'hD5; mem['h0E12]=8'h16; mem['h0E13]=8'hCE;
    mem['h0E14]=8'h44; mem['h0E15]=8'h96; mem['h0E16]=8'h02; mem['h0E17]=8'h36;
    mem['h0E18]=8'h82; mem['h0E19]=8'h2E; mem['h0E1A]=8'h16; mem['h0E1B]=8'hCF;
    mem['h0E1C]=8'h08; mem['h0E1D]=8'h36; mem['h0E1E]=8'hBE; mem['h0E1F]=8'hF9;
    mem['h0E20]=8'h46; mem['h0E21]=8'hAD; mem['h0E22]=8'h02; mem['h0E23]=8'h36;
    mem['h0E24]=8'hD0; mem['h0E25]=8'h2E; mem['h0E26]=8'h01; mem['h0E27]=8'h46;
    mem['h0E28]=8'h0A; mem['h0E29]=8'h0B; mem['h0E2A]=8'hC4; mem['h0E2B]=8'hA0;
    mem['h0E2C]=8'h48; mem['h0E2D]=8'h42; mem['h0E2E]=8'h0E; mem['h0E2F]=8'h36;
    mem['h0E30]=8'h0B; mem['h0E31]=8'h2E; mem['h0E32]=8'h17; mem['h0E33]=8'h46;
    mem['h0E34]=8'h0A; mem['h0E35]=8'h0B; mem['h0E36]=8'hC4; mem['h0E37]=8'hA0;
    mem['h0E38]=8'h48; mem['h0E39]=8'h42; mem['h0E3A]=8'h0E; mem['h0E3B]=8'h06;
    mem['h0E3C]=8'hC9; mem['h0E3D]=8'h16; mem['h0E3E]=8'hC6; mem['h0E3F]=8'h44;
    mem['h0E40]=8'h96; mem['h0E41]=8'h02; mem['h0E42]=8'h36; mem['h0E43]=8'hBF;
    mem['h0E44]=8'h2E; mem['h0E45]=8'h16; mem['h0E46]=8'h21; mem['h0E47]=8'hFC;
    mem['h0E48]=8'h46; mem['h0E49]=8'h94; mem['h0E4A]=8'h03; mem['h0E4B]=8'h36;
    mem['h0E4C]=8'h56; mem['h0E4D]=8'h2E; mem['h0E4E]=8'h01; mem['h0E4F]=8'hC7;
    mem['h0E50]=8'hA0; mem['h0E51]=8'h68; mem['h0E52]=8'h4E; mem['h0E53]=8'h0B;
    mem['h0E54]=8'h36; mem['h0E55]=8'hBF; mem['h0E56]=8'h2E; mem['h0E57]=8'h16;
    mem['h0E58]=8'hC7; mem['h0E59]=8'h04; mem['h0E5A]=8'h05; mem['h0E5B]=8'h36;
    mem['h0E5C]=8'h82; mem['h0E5D]=8'hF8; mem['h0E5E]=8'hC8; mem['h0E5F]=8'h08;
    mem['h0E60]=8'h36; mem['h0E61]=8'h84; mem['h0E62]=8'hF9; mem['h0E63]=8'h36;
    mem['h0E64]=8'h84; mem['h0E65]=8'h46; mem['h0E66]=8'hA0; mem['h0E67]=8'h02;
    mem['h0E68]=8'h48; mem['h0E69]=8'h76; mem['h0E6A]=8'h0E; mem['h0E6B]=8'h36;
    mem['h0E6C]=8'h84; mem['h0E6D]=8'h46; mem['h0E6E]=8'h03; mem['h0E6F]=8'h03;
    mem['h0E70]=8'h48; mem['h0E71]=8'h63; mem['h0E72]=8'h0E; mem['h0E73]=8'h44;
    mem['h0E74]=8'h3B; mem['h0E75]=8'h0E; mem['h0E76]=8'h3C; mem['h0E77]=8'hB0;
    mem['h0E78]=8'h70; mem['h0E79]=8'h80; mem['h0E7A]=8'h0E; mem['h0E7B]=8'h3C;
    mem['h0E7C]=8'hBA; mem['h0E7D]=8'h70; mem['h0E7E]=8'h7C; mem['h0E7F]=8'h0D;
    mem['h0E80]=8'h36; mem['h0E81]=8'h00; mem['h0E82]=8'hC7; mem['h0E83]=8'h36;
    mem['h0E84]=8'h84; mem['h0E85]=8'h97; mem['h0E86]=8'hC8; mem['h0E87]=8'h08;
    mem['h0E88]=8'hD7; mem['h0E89]=8'h36; mem['h0E8A]=8'h00; mem['h0E8B]=8'hF9;
    mem['h0E8C]=8'hF2; mem['h0E8D]=8'h1E; mem['h0E8E]=8'h16; mem['h0E8F]=8'h26;
    mem['h0E90]=8'h01; mem['h0E91]=8'h46; mem['h0E92]=8'h0B; mem['h0E93]=8'h11;
    mem['h0E94]=8'h36; mem['h0E95]=8'h82; mem['h0E96]=8'h3E; mem['h0E97]=8'h01;
    mem['h0E98]=8'h46; mem['h0E99]=8'h37; mem['h0E9A]=8'h02; mem['h0E9B]=8'h44;
    mem['h0E9C]=8'h89; mem['h0E9D]=8'h0B; mem['h0E9E]=8'h36; mem['h0E9F]=8'hE0;
    mem['h0EA0]=8'h2E; mem['h0EA1]=8'h16; mem['h0EA2]=8'hDF; mem['h0EA3]=8'h18;
    mem['h0EA4]=8'h19; mem['h0EA5]=8'h68; mem['h0EA6]=8'hAD; mem['h0EA7]=8'h0E;
    mem['h0EA8]=8'h36; mem['h0EA9]=8'hF0; mem['h0EAA]=8'hDF; mem['h0EAB]=8'h30;
    mem['h0EAC]=8'hE7; mem['h0EAD]=8'h36; mem['h0EAE]=8'h3B; mem['h0EAF]=8'h2E;
    mem['h0EB0]=8'h17; mem['h0EB1]=8'hC7; mem['h0EB2]=8'h04; mem['h0EB3]=8'h02;
    mem['h0EB4]=8'h3C; mem['h0EB5]=8'h11; mem['h0EB6]=8'h50; mem['h0EB7]=8'hE7;
    mem['h0EB8]=8'h0E; mem['h0EB9]=8'hF8; mem['h0EBA]=8'h36; mem['h0EBB]=8'h3E;
    mem['h0EBC]=8'h86; mem['h0EBD]=8'hF0; mem['h0EBE]=8'hFB; mem['h0EBF]=8'h30;
    mem['h0EC0]=8'hFC; mem['h0EC1]=8'h44; mem['h0EC2]=8'h7C; mem['h0EC3]=8'h0D;
    mem['h0EC4]=8'h36; mem['h0EC5]=8'h3B; mem['h0EC6]=8'h2E; mem['h0EC7]=8'h17;
    mem['h0EC8]=8'hC7; mem['h0EC9]=8'h14; mem['h0ECA]=8'h02; mem['h0ECB]=8'h70;
    mem['h0ECC]=8'hEE; mem['h0ECD]=8'h0E; mem['h0ECE]=8'hF8; mem['h0ECF]=8'h04;
    mem['h0ED0]=8'h02; mem['h0ED1]=8'h36; mem['h0ED2]=8'h3E; mem['h0ED3]=8'h86;
    mem['h0ED4]=8'hF0; mem['h0ED5]=8'hDF; mem['h0ED6]=8'h18; mem['h0ED7]=8'h19;
    mem['h0ED8]=8'h68; mem['h0ED9]=8'hB6; mem['h0EDA]=8'h08; mem['h0EDB]=8'h30;
    mem['h0EDC]=8'hE7; mem['h0EDD]=8'h36; mem['h0EDE]=8'hF0; mem['h0EDF]=8'h2E;
    mem['h0EE0]=8'h16; mem['h0EE1]=8'hFB; mem['h0EE2]=8'h30; mem['h0EE3]=8'hFC;
    mem['h0EE4]=8'h44; mem['h0EE5]=8'h4E; mem['h0EE6]=8'h0B; mem['h0EE7]=8'h06;
    mem['h0EE8]=8'hC7; mem['h0EE9]=8'h16; mem['h0EEA]=8'hD3; mem['h0EEB]=8'h44;
    mem['h0EEC]=8'h96; mem['h0EED]=8'h02; mem['h0EEE]=8'h06; mem['h0EEF]=8'hD2;
    mem['h0EF0]=8'h16; mem['h0EF1]=8'hD4; mem['h0EF2]=8'h44; mem['h0EF3]=8'h96;
    mem['h0EF4]=8'h02; mem['h0EF5]=8'h46; mem['h0EF6]=8'hAD; mem['h0EF7]=8'h02;
    mem['h0EF8]=8'h36; mem['h0EF9]=8'h82; mem['h0EFA]=8'hCF; mem['h0EFB]=8'h08;
    mem['h0EFC]=8'h36; mem['h0EFD]=8'h83; mem['h0EFE]=8'hF9; mem['h0EFF]=8'h36;
    mem['h0F00]=8'h83; mem['h0F01]=8'h46; mem['h0F02]=8'hA0; mem['h0F03]=8'h02;
    mem['h0F04]=8'h68; mem['h0F05]=8'h22; mem['h0F06]=8'h0F; mem['h0F07]=8'h3C;
    mem['h0F08]=8'hAC; mem['h0F09]=8'h68; mem['h0F0A]=8'h33; mem['h0F0B]=8'h0F;
    mem['h0F0C]=8'h3C; mem['h0F0D]=8'hA8; mem['h0F0E]=8'h48; mem['h0F0F]=8'h1F;
    mem['h0F10]=8'h0F; mem['h0F11]=8'h46; mem['h0F12]=8'h70; mem['h0F13]=8'h2D;
    mem['h0F14]=8'h36; mem['h0F15]=8'h86; mem['h0F16]=8'h2E; mem['h0F17]=8'h16;
    mem['h0F18]=8'hCF; mem['h0F19]=8'h36; mem['h0F1A]=8'h83; mem['h0F1B]=8'hF9;
    mem['h0F1C]=8'h44; mem['h0F1D]=8'h22; mem['h0F1E]=8'h0F; mem['h0F1F]=8'h46;
    mem['h0F20]=8'hC8; mem['h0F21]=8'h02; mem['h0F22]=8'h36; mem['h0F23]=8'h83;
    mem['h0F24]=8'h46; mem['h0F25]=8'h03; mem['h0F26]=8'h03; mem['h0F27]=8'h48;
    mem['h0F28]=8'hFF; mem['h0F29]=8'h0E; mem['h0F2A]=8'h46; mem['h0F2B]=8'h44;
    mem['h0F2C]=8'h0F; mem['h0F2D]=8'h46; mem['h0F2E]=8'h2D; mem['h0F2F]=8'h08;
    mem['h0F30]=8'h44; mem['h0F31]=8'h4E; mem['h0F32]=8'h0B; mem['h0F33]=8'h46;
    mem['h0F34]=8'h44; mem['h0F35]=8'h0F; mem['h0F36]=8'h46; mem['h0F37]=8'h2D;
    mem['h0F38]=8'h08; mem['h0F39]=8'h2E; mem['h0F3A]=8'h16; mem['h0F3B]=8'h36;
    mem['h0F3C]=8'h83; mem['h0F3D]=8'hCF; mem['h0F3E]=8'h36; mem['h0F3F]=8'h82;
    mem['h0F40]=8'hF9; mem['h0F41]=8'h44; mem['h0F42]=8'hF5; mem['h0F43]=8'h0E;
    mem['h0F44]=8'h36; mem['h0F45]=8'h50; mem['h0F46]=8'hC7; mem['h0F47]=8'h86;
    mem['h0F48]=8'hF0; mem['h0F49]=8'hC7; mem['h0F4A]=8'h3C; mem['h0F4B]=8'hA4;
    mem['h0F4C]=8'h48; mem['h0F4D]=8'h60; mem['h0F4E]=8'h0F; mem['h0F4F]=8'h36;
    mem['h0F50]=8'h50; mem['h0F51]=8'hCF; mem['h0F52]=8'h09; mem['h0F53]=8'hF9;
    mem['h0F54]=8'h46; mem['h0F55]=8'h6F; mem['h0F56]=8'h0F; mem['h0F57]=8'h46;
    mem['h0F58]=8'h91; mem['h0F59]=8'h03; mem['h0F5A]=8'h36; mem['h0F5B]=8'h54;
    mem['h0F5C]=8'hF8; mem['h0F5D]=8'h44; mem['h0F5E]=8'h34; mem['h0F5F]=8'h10;
    mem['h0F60]=8'h36; mem['h0F61]=8'h64; mem['h0F62]=8'h2E; mem['h0F63]=8'h16;
    mem['h0F64]=8'h06; mem['h0F65]=8'hBF; mem['h0F66]=8'h46; mem['h0F67]=8'h82;
    mem['h0F68]=8'h03; mem['h0F69]=8'h46; mem['h0F6A]=8'h0C; mem['h0F6B]=8'h03;
    mem['h0F6C]=8'h44; mem['h0F6D]=8'h24; mem['h0F6E]=8'h13; mem['h0F6F]=8'h2E;
    mem['h0F70]=8'h01; mem['h0F71]=8'h44; mem['h0F72]=8'hA7; mem['h0F73]=8'h06;
    mem['h0F74]=8'h36; mem['h0F75]=8'h64; mem['h0F76]=8'h2E; mem['h0F77]=8'h16;
    mem['h0F78]=8'h3E; mem['h0F79]=8'h00; mem['h0F7A]=8'h36; mem['h0F7B]=8'h66;
    mem['h0F7C]=8'h3E; mem['h0F7D]=8'h00; mem['h0F7E]=8'h36; mem['h0F7F]=8'h85;
    mem['h0F80]=8'h2E; mem['h0F81]=8'h17; mem['h0F82]=8'hCF; mem['h0F83]=8'h08;
    mem['h0F84]=8'hF9; mem['h0F85]=8'h36; mem['h0F86]=8'hF0; mem['h0F87]=8'h2E;
    mem['h0F88]=8'h16; mem['h0F89]=8'hDF; mem['h0F8A]=8'h30; mem['h0F8B]=8'hE7;
    mem['h0F8C]=8'hC1; mem['h0F8D]=8'h02; mem['h0F8E]=8'h02; mem['h0F8F]=8'h04;
    mem['h0F90]=8'h5C; mem['h0F91]=8'hF0; mem['h0F92]=8'h2E; mem['h0F93]=8'h17;
    mem['h0F94]=8'hFB; mem['h0F95]=8'h30; mem['h0F96]=8'hFC; mem['h0F97]=8'h36;
    mem['h0F98]=8'hD5; mem['h0F99]=8'h2E; mem['h0F9A]=8'h01; mem['h0F9B]=8'h46;
    mem['h0F9C]=8'h0A; mem['h0F9D]=8'h0B; mem['h0F9E]=8'hC4; mem['h0F9F]=8'hA0;
    mem['h0FA0]=8'h48; mem['h0FA1]=8'hAA; mem['h0FA2]=8'h0F; mem['h0FA3]=8'h06;
    mem['h0FA4]=8'hC6; mem['h0FA5]=8'h16; mem['h0FA6]=8'hC5; mem['h0FA7]=8'h44;
    mem['h0FA8]=8'h96; mem['h0FA9]=8'h02; mem['h0FAA]=8'h36; mem['h0FAB]=8'h82;
    mem['h0FAC]=8'h2E; mem['h0FAD]=8'h16; mem['h0FAE]=8'hCF; mem['h0FAF]=8'h08;
    mem['h0FB0]=8'h36; mem['h0FB1]=8'h84; mem['h0FB2]=8'hF9; mem['h0FB3]=8'h36;
    mem['h0FB4]=8'h83; mem['h0FB5]=8'hFC; mem['h0FB6]=8'h36; mem['h0FB7]=8'h84;
    mem['h0FB8]=8'h46; mem['h0FB9]=8'hA0; mem['h0FBA]=8'h02; mem['h0FBB]=8'h68;
    mem['h0FBC]=8'hC8; mem['h0FBD]=8'h0F; mem['h0FBE]=8'h3C; mem['h0FBF]=8'hBD;
    mem['h0FC0]=8'h68; mem['h0FC1]=8'hD3; mem['h0FC2]=8'h0F; mem['h0FC3]=8'h36;
    mem['h0FC4]=8'h64; mem['h0FC5]=8'h46; mem['h0FC6]=8'hCC; mem['h0FC7]=8'h02;
    mem['h0FC8]=8'h36; mem['h0FC9]=8'h84; mem['h0FCA]=8'h46; mem['h0FCB]=8'h03;
    mem['h0FCC]=8'h03; mem['h0FCD]=8'h48; mem['h0FCE]=8'hB6; mem['h0FCF]=8'h0F;
    mem['h0FD0]=8'h44; mem['h0FD1]=8'hA3; mem['h0FD2]=8'h0F; mem['h0FD3]=8'h36;
    mem['h0FD4]=8'h84; mem['h0FD5]=8'hCF; mem['h0FD6]=8'h08; mem['h0FD7]=8'h36;
    mem['h0FD8]=8'hBE; mem['h0FD9]=8'hF9; mem['h0FDA]=8'h36; mem['h0FDB]=8'h83;
    mem['h0FDC]=8'hCF; mem['h0FDD]=8'h09; mem['h0FDE]=8'h36; mem['h0FDF]=8'hBF;
    mem['h0FE0]=8'hF9; mem['h0FE1]=8'h46; mem['h0FE2]=8'h94; mem['h0FE3]=8'h03;
    mem['h0FE4]=8'h46; mem['h0FE5]=8'hAA; mem['h0FE6]=8'h08; mem['h0FE7]=8'h36;
    mem['h0FE8]=8'h64; mem['h0FE9]=8'h2E; mem['h0FEA]=8'h16; mem['h0FEB]=8'hC7;
    mem['h0FEC]=8'h3C; mem['h0FED]=8'h01; mem['h0FEE]=8'h48; mem['h0FEF]=8'hA6;
    mem['h0FF0]=8'h19; mem['h0FF1]=8'h36; mem['h0FF2]=8'h66; mem['h0FF3]=8'h3E;
    mem['h0FF4]=8'h00; mem['h0FF5]=8'h44; mem['h0FF6]=8'hA6; mem['h0FF7]=8'h19;
    mem['h0FF8]=8'hFF; mem['h0FF9]=8'hFF; mem['h0FFA]=8'hFF; mem['h0FFB]=8'hFF;
    mem['h0FFC]=8'hFF; mem['h0FFD]=8'hFF; mem['h0FFE]=8'hFF; mem['h0FFF]=8'hFF;
    mem['h1000]=8'h36; mem['h1001]=8'h56; mem['h1002]=8'h2E; mem['h1003]=8'h01;
    mem['h1004]=8'hC7; mem['h1005]=8'h36; mem['h1006]=8'h40; mem['h1007]=8'hF8;
    mem['h1008]=8'hA0; mem['h1009]=8'h72; mem['h100A]=8'h82; mem['h100B]=8'h10;
    mem['h100C]=8'h36; mem['h100D]=8'h57; mem['h100E]=8'h06; mem['h100F]=8'h17;
    mem['h1010]=8'hCF; mem['h1011]=8'h08; mem['h1012]=8'h09; mem['h1013]=8'h70;
    mem['h1014]=8'h29; mem['h1015]=8'h10; mem['h1016]=8'h91; mem['h1017]=8'h70;
    mem['h1018]=8'hF6; mem['h1019]=8'h0A; mem['h101A]=8'hD0; mem['h101B]=8'h36;
    mem['h101C]=8'h56; mem['h101D]=8'h0E; mem['h101E]=8'h03; mem['h101F]=8'h46;
    mem['h1020]=8'h89; mem['h1021]=8'h12; mem['h1022]=8'h11; mem['h1023]=8'h48;
    mem['h1024]=8'h1B; mem['h1025]=8'h10; mem['h1026]=8'h44; mem['h1027]=8'h7D;
    mem['h1028]=8'h10; mem['h1029]=8'h36; mem['h102A]=8'h56; mem['h102B]=8'hA8;
    mem['h102C]=8'hF8; mem['h102D]=8'h31; mem['h102E]=8'hF8; mem['h102F]=8'h31;
    mem['h1030]=8'hF8; mem['h1031]=8'h31; mem['h1032]=8'hF8; mem['h1033]=8'h07;
    mem['h1034]=8'h0E; mem['h1035]=8'h17; mem['h1036]=8'hC1; mem['h1037]=8'h2E;
    mem['h1038]=8'h01; mem['h1039]=8'h36; mem['h103A]=8'h57; mem['h103B]=8'hA0;
    mem['h103C]=8'h68; mem['h103D]=8'h40; mem['h103E]=8'h10; mem['h103F]=8'hF9;
    mem['h1040]=8'h31; mem['h1041]=8'hC7; mem['h1042]=8'h36; mem['h1043]=8'h40;
    mem['h1044]=8'hF8; mem['h1045]=8'hA0; mem['h1046]=8'h50; mem['h1047]=8'h50;
    mem['h1048]=8'h10; mem['h1049]=8'h0E; mem['h104A]=8'h04; mem['h104B]=8'h36;
    mem['h104C]=8'h53; mem['h104D]=8'h46; mem['h104E]=8'h68; mem['h104F]=8'h12;
    mem['h1050]=8'h36; mem['h1051]=8'h56; mem['h1052]=8'h0E; mem['h1053]=8'h04;
    mem['h1054]=8'hC7; mem['h1055]=8'hA0; mem['h1056]=8'h48; mem['h1057]=8'h63;
    mem['h1058]=8'h10; mem['h1059]=8'h31; mem['h105A]=8'h09; mem['h105B]=8'h48;
    mem['h105C]=8'h54; mem['h105D]=8'h10; mem['h105E]=8'h36; mem['h105F]=8'h57;
    mem['h1060]=8'hA8; mem['h1061]=8'hF8; mem['h1062]=8'h07; mem['h1063]=8'h36;
    mem['h1064]=8'h53; mem['h1065]=8'h0E; mem['h1066]=8'h04; mem['h1067]=8'h46;
    mem['h1068]=8'h7F; mem['h1069]=8'h12; mem['h106A]=8'hC7; mem['h106B]=8'hA0;
    mem['h106C]=8'h70; mem['h106D]=8'h76; mem['h106E]=8'h10; mem['h106F]=8'h30;
    mem['h1070]=8'hCF; mem['h1071]=8'h09; mem['h1072]=8'hF9; mem['h1073]=8'h44;
    mem['h1074]=8'h63; mem['h1075]=8'h10; mem['h1076]=8'h36; mem['h1077]=8'h56;
    mem['h1078]=8'h0E; mem['h1079]=8'h03; mem['h107A]=8'h46; mem['h107B]=8'h89;
    mem['h107C]=8'h12; mem['h107D]=8'h36; mem['h107E]=8'h40; mem['h107F]=8'hC7;
    mem['h1080]=8'hA0; mem['h1081]=8'h13; mem['h1082]=8'h36; mem['h1083]=8'h54;
    mem['h1084]=8'h0E; mem['h1085]=8'h03; mem['h1086]=8'h44; mem['h1087]=8'h68;
    mem['h1088]=8'h12; mem['h1089]=8'h36; mem['h108A]=8'h56; mem['h108B]=8'h2E;
    mem['h108C]=8'h01; mem['h108D]=8'hC7; mem['h108E]=8'hA0; mem['h108F]=8'h48;
    mem['h1090]=8'h9D; mem['h1091]=8'h10; mem['h1092]=8'h36; mem['h1093]=8'h54;
    mem['h1094]=8'hDD; mem['h1095]=8'hE6; mem['h1096]=8'h36; mem['h1097]=8'h5C;
    mem['h1098]=8'h0E; mem['h1099]=8'h04; mem['h109A]=8'h44; mem['h109B]=8'h0B;
    mem['h109C]=8'h11; mem['h109D]=8'h36; mem['h109E]=8'h5E; mem['h109F]=8'hC7;
    mem['h10A0]=8'hA0; mem['h10A1]=8'h2B; mem['h10A2]=8'h36; mem['h10A3]=8'h57;
    mem['h10A4]=8'hC7; mem['h10A5]=8'h36; mem['h10A6]=8'h5F; mem['h10A7]=8'hBF;
    mem['h10A8]=8'h68; mem['h10A9]=8'hE1; mem['h10AA]=8'h10; mem['h10AB]=8'hC8;
    mem['h10AC]=8'hC7; mem['h10AD]=8'h99; mem['h10AE]=8'h50; mem['h10AF]=8'hB4;
    mem['h10B0]=8'h10; mem['h10B1]=8'hC8; mem['h10B2]=8'hA8; mem['h10B3]=8'h99;
    mem['h10B4]=8'h3C; mem['h10B5]=8'h18; mem['h10B6]=8'h70; mem['h10B7]=8'hC3;
    mem['h10B8]=8'h10; mem['h10B9]=8'hC7; mem['h10BA]=8'h36; mem['h10BB]=8'h57;
    mem['h10BC]=8'h97; mem['h10BD]=8'h33; mem['h10BE]=8'h36; mem['h10BF]=8'h54;
    mem['h10C0]=8'h44; mem['h10C1]=8'h92; mem['h10C2]=8'h10; mem['h10C3]=8'hC7;
    mem['h10C4]=8'h36; mem['h10C5]=8'h57; mem['h10C6]=8'h97; mem['h10C7]=8'h70;
    mem['h10C8]=8'hD7; mem['h10C9]=8'h10; mem['h10CA]=8'hD0; mem['h10CB]=8'h36;
    mem['h10CC]=8'h57; mem['h10CD]=8'h46; mem['h10CE]=8'hFC; mem['h10CF]=8'h10;
    mem['h10D0]=8'h11; mem['h10D1]=8'h48; mem['h10D2]=8'hCB; mem['h10D3]=8'h10;
    mem['h10D4]=8'h44; mem['h10D5]=8'hE1; mem['h10D6]=8'h10; mem['h10D7]=8'hD0;
    mem['h10D8]=8'h36; mem['h10D9]=8'h5F; mem['h10DA]=8'h46; mem['h10DB]=8'hFC;
    mem['h10DC]=8'h10; mem['h10DD]=8'h10; mem['h10DE]=8'h48; mem['h10DF]=8'hD8;
    mem['h10E0]=8'h10; mem['h10E1]=8'h46; mem['h10E2]=8'h00; mem['h10E3]=8'h18;
    mem['h10E4]=8'hC0; mem['h10E5]=8'h36; mem['h10E6]=8'h57; mem['h10E7]=8'h46;
    mem['h10E8]=8'hFC; mem['h10E9]=8'h10; mem['h10EA]=8'h36; mem['h10EB]=8'h5F;
    mem['h10EC]=8'h46; mem['h10ED]=8'hFC; mem['h10EE]=8'h10; mem['h10EF]=8'hDD;
    mem['h10F0]=8'h26; mem['h10F1]=8'h53; mem['h10F2]=8'h0E; mem['h10F3]=8'h04;
    mem['h10F4]=8'h46; mem['h10F5]=8'h57; mem['h10F6]=8'h12; mem['h10F7]=8'h0E;
    mem['h10F8]=8'h00; mem['h10F9]=8'h44; mem['h10FA]=8'h36; mem['h10FB]=8'h10;
    mem['h10FC]=8'hCF; mem['h10FD]=8'h08; mem['h10FE]=8'hF9; mem['h10FF]=8'h31;
    mem['h1100]=8'h0E; mem['h1101]=8'h04; mem['h1102]=8'hC7; mem['h1103]=8'hA0;
    mem['h1104]=8'h50; mem['h1105]=8'h89; mem['h1106]=8'h12; mem['h1107]=8'h12;
    mem['h1108]=8'h44; mem['h1109]=8'h8A; mem['h110A]=8'h12; mem['h110B]=8'hC7;
    mem['h110C]=8'h30; mem['h110D]=8'h46; mem['h110E]=8'hEE; mem['h110F]=8'h12;
    mem['h1110]=8'hF8; mem['h1111]=8'h30; mem['h1112]=8'h46; mem['h1113]=8'hEE;
    mem['h1114]=8'h12; mem['h1115]=8'h09; mem['h1116]=8'h2B; mem['h1117]=8'h44;
    mem['h1118]=8'h0B; mem['h1119]=8'h11; mem['h111A]=8'h36; mem['h111B]=8'h54;
    mem['h111C]=8'h2E; mem['h111D]=8'h01; mem['h111E]=8'h0E; mem['h111F]=8'h03;
    mem['h1120]=8'h46; mem['h1121]=8'h68; mem['h1122]=8'h12; mem['h1123]=8'h44;
    mem['h1124]=8'h89; mem['h1125]=8'h10; mem['h1126]=8'h46; mem['h1127]=8'h76;
    mem['h1128]=8'h11; mem['h1129]=8'h36; mem['h112A]=8'h5F; mem['h112B]=8'hC7;
    mem['h112C]=8'h36; mem['h112D]=8'h57; mem['h112E]=8'h87; mem['h112F]=8'h04;
    mem['h1130]=8'h01; mem['h1131]=8'hF8; mem['h1132]=8'h36; mem['h1133]=8'h42;
    mem['h1134]=8'h3E; mem['h1135]=8'h17; mem['h1136]=8'h36; mem['h1137]=8'h56;
    mem['h1138]=8'h0E; mem['h1139]=8'h03; mem['h113A]=8'h46; mem['h113B]=8'h89;
    mem['h113C]=8'h12; mem['h113D]=8'h62; mem['h113E]=8'hB8; mem['h113F]=8'h11;
    mem['h1140]=8'h36; mem['h1141]=8'h66; mem['h1142]=8'h0E; mem['h1143]=8'h06;
    mem['h1144]=8'h46; mem['h1145]=8'h89; mem['h1146]=8'h12; mem['h1147]=8'h36;
    mem['h1148]=8'h42; mem['h1149]=8'hD7; mem['h114A]=8'h11; mem['h114B]=8'hFA;
    mem['h114C]=8'h48; mem['h114D]=8'h36; mem['h114E]=8'h11; mem['h114F]=8'h36;
    mem['h1150]=8'h66; mem['h1151]=8'h0E; mem['h1152]=8'h06; mem['h1153]=8'h46;
    mem['h1154]=8'h89; mem['h1155]=8'h12; mem['h1156]=8'h36; mem['h1157]=8'h63;
    mem['h1158]=8'hC7; mem['h1159]=8'h12; mem['h115A]=8'hA0; mem['h115B]=8'h72;
    mem['h115C]=8'hC2; mem['h115D]=8'h11; mem['h115E]=8'h36; mem['h115F]=8'h53;
    mem['h1160]=8'hE6; mem['h1161]=8'hDD; mem['h1162]=8'h36; mem['h1163]=8'h63;
    mem['h1164]=8'h0E; mem['h1165]=8'h04; mem['h1166]=8'h46; mem['h1167]=8'h0B;
    mem['h1168]=8'h11; mem['h1169]=8'h0E; mem['h116A]=8'h00; mem['h116B]=8'h46;
    mem['h116C]=8'h36; mem['h116D]=8'h10; mem['h116E]=8'h36; mem['h116F]=8'h41;
    mem['h1170]=8'hC7; mem['h1171]=8'hA0; mem['h1172]=8'h0B; mem['h1173]=8'h44;
    mem['h1174]=8'h82; mem['h1175]=8'h10; mem['h1176]=8'h36; mem['h1177]=8'h60;
    mem['h1178]=8'h2E; mem['h1179]=8'h01; mem['h117A]=8'h0E; mem['h117B]=8'h08;
    mem['h117C]=8'hA8; mem['h117D]=8'hF8; mem['h117E]=8'h30; mem['h117F]=8'h09;
    mem['h1180]=8'h48; mem['h1181]=8'h7D; mem['h1182]=8'h11; mem['h1183]=8'h0E;
    mem['h1184]=8'h04; mem['h1185]=8'h36; mem['h1186]=8'h58; mem['h1187]=8'hF8;
    mem['h1188]=8'h30; mem['h1189]=8'h09; mem['h118A]=8'h48; mem['h118B]=8'h87;
    mem['h118C]=8'h11; mem['h118D]=8'h36; mem['h118E]=8'h41; mem['h118F]=8'h3E;
    mem['h1190]=8'h01; mem['h1191]=8'h36; mem['h1192]=8'h56; mem['h1193]=8'hC7;
    mem['h1194]=8'hA0; mem['h1195]=8'h70; mem['h1196]=8'hA9; mem['h1197]=8'h11;
    mem['h1198]=8'h36; mem['h1199]=8'h5E; mem['h119A]=8'hC7; mem['h119B]=8'hA0;
    mem['h119C]=8'h13; mem['h119D]=8'h36; mem['h119E]=8'h41; mem['h119F]=8'hD7;
    mem['h11A0]=8'h11; mem['h11A1]=8'hFA; mem['h11A2]=8'h36; mem['h11A3]=8'h5C;
    mem['h11A4]=8'h0E; mem['h11A5]=8'h03; mem['h11A6]=8'h44; mem['h11A7]=8'h68;
    mem['h11A8]=8'h12; mem['h11A9]=8'h36; mem['h11AA]=8'h41; mem['h11AB]=8'hD7;
    mem['h11AC]=8'h11; mem['h11AD]=8'hFA; mem['h11AE]=8'h36; mem['h11AF]=8'h54;
    mem['h11B0]=8'h0E; mem['h11B1]=8'h03; mem['h11B2]=8'h46; mem['h11B3]=8'h68;
    mem['h11B4]=8'h12; mem['h11B5]=8'h44; mem['h11B6]=8'h98; mem['h11B7]=8'h11;
    mem['h11B8]=8'h26; mem['h11B9]=8'h61; mem['h11BA]=8'hDD; mem['h11BB]=8'h36;
    mem['h11BC]=8'h59; mem['h11BD]=8'h0E; mem['h11BE]=8'h06; mem['h11BF]=8'h44;
    mem['h11C0]=8'h57; mem['h11C1]=8'h12; mem['h11C2]=8'h0E; mem['h11C3]=8'h03;
    mem['h11C4]=8'h06; mem['h11C5]=8'h40; mem['h11C6]=8'h87; mem['h11C7]=8'hF8;
    mem['h11C8]=8'h30; mem['h11C9]=8'h06; mem['h11CA]=8'h00; mem['h11CB]=8'h8F;
    mem['h11CC]=8'h09; mem['h11CD]=8'h48; mem['h11CE]=8'hC7; mem['h11CF]=8'h11;
    mem['h11D0]=8'hF8; mem['h11D1]=8'h07; mem['h11D2]=8'h46; mem['h11D3]=8'h76;
    mem['h11D4]=8'h11; mem['h11D5]=8'h36; mem['h11D6]=8'h56; mem['h11D7]=8'hC7;
    mem['h11D8]=8'hA0; mem['h11D9]=8'h68; mem['h11DA]=8'hEF; mem['h11DB]=8'h0A;
    mem['h11DC]=8'h36; mem['h11DD]=8'h5F; mem['h11DE]=8'hC7; mem['h11DF]=8'h36;
    mem['h11E0]=8'h57; mem['h11E1]=8'h97; mem['h11E2]=8'h04; mem['h11E3]=8'h01;
    mem['h11E4]=8'hF8; mem['h11E5]=8'h36; mem['h11E6]=8'h42; mem['h11E7]=8'h3E;
    mem['h11E8]=8'h17; mem['h11E9]=8'h46; mem['h11EA]=8'h41; mem['h11EB]=8'h12;
    mem['h11EC]=8'h70; mem['h11ED]=8'hFE; mem['h11EE]=8'h11; mem['h11EF]=8'h26;
    mem['h11F0]=8'h5C; mem['h11F1]=8'h36; mem['h11F2]=8'h59; mem['h11F3]=8'h0E;
    mem['h11F4]=8'h03; mem['h11F5]=8'h46; mem['h11F6]=8'h0B; mem['h11F7]=8'h11;
    mem['h11F8]=8'h06; mem['h11F9]=8'h01; mem['h11FA]=8'h1A; mem['h11FB]=8'h44;
    mem['h11FC]=8'hFF; mem['h11FD]=8'h11; mem['h11FE]=8'hA8; mem['h11FF]=8'h36;
    mem['h1200]=8'h64; mem['h1201]=8'h0E; mem['h1202]=8'h03; mem['h1203]=8'h46;
    mem['h1204]=8'h80; mem['h1205]=8'h12; mem['h1206]=8'h36; mem['h1207]=8'h5C;
    mem['h1208]=8'h0E; mem['h1209]=8'h03; mem['h120A]=8'h46; mem['h120B]=8'h7F;
    mem['h120C]=8'h12; mem['h120D]=8'h36; mem['h120E]=8'h42; mem['h120F]=8'hD7;
    mem['h1210]=8'h11; mem['h1211]=8'hFA; mem['h1212]=8'h48; mem['h1213]=8'hE9;
    mem['h1214]=8'h11; mem['h1215]=8'h46; mem['h1216]=8'h41; mem['h1217]=8'h12;
    mem['h1218]=8'h70; mem['h1219]=8'h38; mem['h121A]=8'h12; mem['h121B]=8'h36;
    mem['h121C]=8'h64; mem['h121D]=8'hC7; mem['h121E]=8'h04; mem['h121F]=8'h01;
    mem['h1220]=8'hF8; mem['h1221]=8'h06; mem['h1222]=8'h00; mem['h1223]=8'h30;
    mem['h1224]=8'h8F; mem['h1225]=8'hF8; mem['h1226]=8'h06; mem['h1227]=8'h00;
    mem['h1228]=8'h30; mem['h1229]=8'h8F; mem['h122A]=8'hF8; mem['h122B]=8'h50;
    mem['h122C]=8'h38; mem['h122D]=8'h12; mem['h122E]=8'h0E; mem['h122F]=8'h03;
    mem['h1230]=8'h46; mem['h1231]=8'h89; mem['h1232]=8'h12; mem['h1233]=8'h36;
    mem['h1234]=8'h57; mem['h1235]=8'hCF; mem['h1236]=8'h08; mem['h1237]=8'hF9;
    mem['h1238]=8'h36; mem['h1239]=8'h63; mem['h123A]=8'h26; mem['h123B]=8'h53;
    mem['h123C]=8'h0E; mem['h123D]=8'h04; mem['h123E]=8'h44; mem['h123F]=8'h66;
    mem['h1240]=8'h11; mem['h1241]=8'h26; mem['h1242]=8'h59; mem['h1243]=8'hDD;
    mem['h1244]=8'h36; mem['h1245]=8'h54; mem['h1246]=8'h0E; mem['h1247]=8'h03;
    mem['h1248]=8'h46; mem['h1249]=8'h0B; mem['h124A]=8'h11; mem['h124B]=8'h26;
    mem['h124C]=8'h59; mem['h124D]=8'h36; mem['h124E]=8'h5C; mem['h124F]=8'h0E;
    mem['h1250]=8'h03; mem['h1251]=8'h46; mem['h1252]=8'h93; mem['h1253]=8'h12;
    mem['h1254]=8'hC7; mem['h1255]=8'hA0; mem['h1256]=8'h07; mem['h1257]=8'hA0;
    mem['h1258]=8'hC7; mem['h1259]=8'h46; mem['h125A]=8'hEE; mem['h125B]=8'h12;
    mem['h125C]=8'h8F; mem['h125D]=8'hF8; mem['h125E]=8'h09; mem['h125F]=8'h2B;
    mem['h1260]=8'h30; mem['h1261]=8'h46; mem['h1262]=8'hEE; mem['h1263]=8'h12;
    mem['h1264]=8'h30; mem['h1265]=8'h44; mem['h1266]=8'h58; mem['h1267]=8'h12;
    mem['h1268]=8'hC7; mem['h1269]=8'h2C; mem['h126A]=8'hFF; mem['h126B]=8'h04;
    mem['h126C]=8'h01; mem['h126D]=8'hF8; mem['h126E]=8'h1A; mem['h126F]=8'hD8;
    mem['h1270]=8'h09; mem['h1271]=8'h2B; mem['h1272]=8'h30; mem['h1273]=8'hC7;
    mem['h1274]=8'h2C; mem['h1275]=8'hFF; mem['h1276]=8'hE0; mem['h1277]=8'hC3;
    mem['h1278]=8'h12; mem['h1279]=8'h06; mem['h127A]=8'h00; mem['h127B]=8'h8C;
    mem['h127C]=8'h44; mem['h127D]=8'h6D; mem['h127E]=8'h12; mem['h127F]=8'hA0;
    mem['h1280]=8'hC7; mem['h1281]=8'h12; mem['h1282]=8'hF8; mem['h1283]=8'h09;
    mem['h1284]=8'h2B; mem['h1285]=8'h30; mem['h1286]=8'h44; mem['h1287]=8'h80;
    mem['h1288]=8'h12; mem['h1289]=8'hA0; mem['h128A]=8'hC7; mem['h128B]=8'h1A;
    mem['h128C]=8'hF8; mem['h128D]=8'h09; mem['h128E]=8'h2B; mem['h128F]=8'h31;
    mem['h1290]=8'h44; mem['h1291]=8'h8A; mem['h1292]=8'h12; mem['h1293]=8'hA0;
    mem['h1294]=8'hC7; mem['h1295]=8'h46; mem['h1296]=8'hEE; mem['h1297]=8'h12;
    mem['h1298]=8'h9F; mem['h1299]=8'hF8; mem['h129A]=8'h09; mem['h129B]=8'h2B;
    mem['h129C]=8'h30; mem['h129D]=8'h46; mem['h129E]=8'hEE; mem['h129F]=8'h12;
    mem['h12A0]=8'h30; mem['h12A1]=8'h44; mem['h12A2]=8'h94; mem['h12A3]=8'h12;
    mem['h12A4]=8'h1E; mem['h12A5]=8'h01; mem['h12A6]=8'h26; mem['h12A7]=8'h54;
    mem['h12A8]=8'h0E; mem['h12A9]=8'h04; mem['h12AA]=8'h44; mem['h12AB]=8'h0B;
    mem['h12AC]=8'h11; mem['h12AD]=8'hE6; mem['h12AE]=8'hDD; mem['h12AF]=8'h36;
    mem['h12B0]=8'h54; mem['h12B1]=8'h2E; mem['h12B2]=8'h01; mem['h12B3]=8'h44;
    mem['h12B4]=8'hBA; mem['h12B5]=8'h12; mem['h12B6]=8'h1E; mem['h12B7]=8'h01;
    mem['h12B8]=8'h26; mem['h12B9]=8'h5C; mem['h12BA]=8'h0E; mem['h12BB]=8'h04;
    mem['h12BC]=8'h44; mem['h12BD]=8'h0B; mem['h12BE]=8'h11; mem['h12BF]=8'h46;
    mem['h12C0]=8'hCF; mem['h12C1]=8'h12; mem['h12C2]=8'h36; mem['h12C3]=8'h54;
    mem['h12C4]=8'h2E; mem['h12C5]=8'h01; mem['h12C6]=8'h46; mem['h12C7]=8'hB6;
    mem['h12C8]=8'h12; mem['h12C9]=8'h46; mem['h12CA]=8'hDF; mem['h12CB]=8'h12;
    mem['h12CC]=8'h44; mem['h12CD]=8'hA4; mem['h12CE]=8'h12; mem['h12CF]=8'hC5;
    mem['h12D0]=8'hCE; mem['h12D1]=8'h36; mem['h12D2]=8'h80; mem['h12D3]=8'h2E;
    mem['h12D4]=8'h01; mem['h12D5]=8'hF8; mem['h12D6]=8'h30; mem['h12D7]=8'hF9;
    mem['h12D8]=8'h30; mem['h12D9]=8'hFB; mem['h12DA]=8'h30; mem['h12DB]=8'hFC;
    mem['h12DC]=8'hE8; mem['h12DD]=8'hF1; mem['h12DE]=8'h07; mem['h12DF]=8'h36;
    mem['h12E0]=8'h80; mem['h12E1]=8'h2E; mem['h12E2]=8'h01; mem['h12E3]=8'hC7;
    mem['h12E4]=8'h30; mem['h12E5]=8'hCF; mem['h12E6]=8'h30; mem['h12E7]=8'hDF;
    mem['h12E8]=8'h30; mem['h12E9]=8'hE7; mem['h12EA]=8'hE8; mem['h12EB]=8'hF1;
    mem['h12EC]=8'hC7; mem['h12ED]=8'h07; mem['h12EE]=8'hD5; mem['h12EF]=8'hEB;
    mem['h12F0]=8'hDA; mem['h12F1]=8'hD6; mem['h12F2]=8'hF4; mem['h12F3]=8'hE2;
    mem['h12F4]=8'h07; mem['h12F5]=8'h2E; mem['h12F6]=8'h01; mem['h12F7]=8'h36;
    mem['h12F8]=8'h90; mem['h12F9]=8'hD7; mem['h12FA]=8'h10; mem['h12FB]=8'h11;
    mem['h12FC]=8'h48; mem['h12FD]=8'h08; mem['h12FE]=8'h13; mem['h12FF]=8'hF4;
    mem['h1300]=8'hEB; mem['h1301]=8'hD7; mem['h1302]=8'h10; mem['h1303]=8'h46;
    mem['h1304]=8'h1E; mem['h1305]=8'h13; mem['h1306]=8'h3E; mem['h1307]=8'h00;
    mem['h1308]=8'h36; mem['h1309]=8'h90; mem['h130A]=8'h2E; mem['h130B]=8'h01;
    mem['h130C]=8'hD7; mem['h130D]=8'h10; mem['h130E]=8'hFA; mem['h130F]=8'hF4;
    mem['h1310]=8'hEB; mem['h1311]=8'h46; mem['h1312]=8'h1E; mem['h1313]=8'h13;
    mem['h1314]=8'hC7; mem['h1315]=8'hA0; mem['h1316]=8'h2E; mem['h1317]=8'h01;
    mem['h1318]=8'h0B; mem['h1319]=8'h36; mem['h131A]=8'h90; mem['h131B]=8'h3E;
    mem['h131C]=8'h00; mem['h131D]=8'h07; mem['h131E]=8'hC6; mem['h131F]=8'h82;
    mem['h1320]=8'hF0; mem['h1321]=8'h03; mem['h1322]=8'h28; mem['h1323]=8'h07;
    mem['h1324]=8'hE6; mem['h1325]=8'hDD; mem['h1326]=8'h2E; mem['h1327]=8'h01;
    mem['h1328]=8'h36; mem['h1329]=8'h68; mem['h132A]=8'hA8; mem['h132B]=8'h0E;
    mem['h132C]=8'h08; mem['h132D]=8'hF8; mem['h132E]=8'h30; mem['h132F]=8'h09;
    mem['h1330]=8'h48; mem['h1331]=8'h2D; mem['h1332]=8'h13; mem['h1333]=8'h36;
    mem['h1334]=8'h43; mem['h1335]=8'h0E; mem['h1336]=8'h04; mem['h1337]=8'hF8;
    mem['h1338]=8'h30; mem['h1339]=8'h09; mem['h133A]=8'h48; mem['h133B]=8'h37;
    mem['h133C]=8'h13; mem['h133D]=8'h46; mem['h133E]=8'hF5; mem['h133F]=8'h12;
    mem['h1340]=8'h3C; mem['h1341]=8'hAB; mem['h1342]=8'h68; mem['h1343]=8'h4D;
    mem['h1344]=8'h13; mem['h1345]=8'h3C; mem['h1346]=8'hAD; mem['h1347]=8'h48;
    mem['h1348]=8'h50; mem['h1349]=8'h13; mem['h134A]=8'h36; mem['h134B]=8'h43;
    mem['h134C]=8'hF8; mem['h134D]=8'h46; mem['h134E]=8'hF5; mem['h134F]=8'h12;
    mem['h1350]=8'h3C; mem['h1351]=8'hAE; mem['h1352]=8'h68; mem['h1353]=8'h81;
    mem['h1354]=8'h13; mem['h1355]=8'h3C; mem['h1356]=8'hC5; mem['h1357]=8'h68;
    mem['h1358]=8'h91; mem['h1359]=8'h13; mem['h135A]=8'h3C; mem['h135B]=8'hA0;
    mem['h135C]=8'h68; mem['h135D]=8'h4D; mem['h135E]=8'h13; mem['h135F]=8'hA0;
    mem['h1360]=8'h68; mem['h1361]=8'hC9; mem['h1362]=8'h13; mem['h1363]=8'h3C;
    mem['h1364]=8'hB0; mem['h1365]=8'h70; mem['h1366]=8'hFD; mem['h1367]=8'h0A;
    mem['h1368]=8'h3C; mem['h1369]=8'hBA; mem['h136A]=8'h50; mem['h136B]=8'hFD;
    mem['h136C]=8'h0A; mem['h136D]=8'h36; mem['h136E]=8'h6E; mem['h136F]=8'hD0;
    mem['h1370]=8'h06; mem['h1371]=8'hF8; mem['h1372]=8'hA7; mem['h1373]=8'h48;
    mem['h1374]=8'h4D; mem['h1375]=8'h13; mem['h1376]=8'h36; mem['h1377]=8'h45;
    mem['h1378]=8'hCF; mem['h1379]=8'h08; mem['h137A]=8'hF9; mem['h137B]=8'h46;
    mem['h137C]=8'h2E; mem['h137D]=8'h14; mem['h137E]=8'h44; mem['h137F]=8'h4D;
    mem['h1380]=8'h13; mem['h1381]=8'hC8; mem['h1382]=8'h36; mem['h1383]=8'h46;
    mem['h1384]=8'hC7; mem['h1385]=8'hA0; mem['h1386]=8'h48; mem['h1387]=8'hFD;
    mem['h1388]=8'h0A; mem['h1389]=8'h36; mem['h138A]=8'h45; mem['h138B]=8'hF8;
    mem['h138C]=8'h30; mem['h138D]=8'hF9; mem['h138E]=8'h44; mem['h138F]=8'h4D;
    mem['h1390]=8'h13; mem['h1391]=8'h46; mem['h1392]=8'hF5; mem['h1393]=8'h12;
    mem['h1394]=8'h3C; mem['h1395]=8'hAB; mem['h1396]=8'h68; mem['h1397]=8'hA1;
    mem['h1398]=8'h13; mem['h1399]=8'h3C; mem['h139A]=8'hAD; mem['h139B]=8'h48;
    mem['h139C]=8'hA4; mem['h139D]=8'h13; mem['h139E]=8'h36; mem['h139F]=8'h44;
    mem['h13A0]=8'hF8; mem['h13A1]=8'h46; mem['h13A2]=8'hF5; mem['h13A3]=8'h12;
    mem['h13A4]=8'hA0; mem['h13A5]=8'h68; mem['h13A6]=8'hC9; mem['h13A7]=8'h13;
    mem['h13A8]=8'h3C; mem['h13A9]=8'hB0; mem['h13AA]=8'h70; mem['h13AB]=8'hFD;
    mem['h13AC]=8'h0A; mem['h13AD]=8'h3C; mem['h13AE]=8'hBA; mem['h13AF]=8'h50;
    mem['h13B0]=8'hFD; mem['h13B1]=8'h0A; mem['h13B2]=8'h24; mem['h13B3]=8'h0F;
    mem['h13B4]=8'hC8; mem['h13B5]=8'h36; mem['h13B6]=8'h6F; mem['h13B7]=8'h06;
    mem['h13B8]=8'h03; mem['h13B9]=8'hBF; mem['h13BA]=8'h70; mem['h13BB]=8'hFD;
    mem['h13BC]=8'h0A; mem['h13BD]=8'hD7; mem['h13BE]=8'hC7; mem['h13BF]=8'hA0;
    mem['h13C0]=8'h12; mem['h13C1]=8'h12; mem['h13C2]=8'h82; mem['h13C3]=8'h12;
    mem['h13C4]=8'h81; mem['h13C5]=8'hF8; mem['h13C6]=8'h44; mem['h13C7]=8'hA1;
    mem['h13C8]=8'h13; mem['h13C9]=8'h36; mem['h13CA]=8'h43; mem['h13CB]=8'hC7;
    mem['h13CC]=8'hA0; mem['h13CD]=8'h68; mem['h13CE]=8'hD7; mem['h13CF]=8'h13;
    mem['h13D0]=8'h36; mem['h13D1]=8'h6C; mem['h13D2]=8'h0E; mem['h13D3]=8'h03;
    mem['h13D4]=8'h46; mem['h13D5]=8'h68; mem['h13D6]=8'h12; mem['h13D7]=8'h36;
    mem['h13D8]=8'h6B; mem['h13D9]=8'hA8; mem['h13DA]=8'hF8; mem['h13DB]=8'hDD;
    mem['h13DC]=8'h26; mem['h13DD]=8'h53; mem['h13DE]=8'h0E; mem['h13DF]=8'h04;
    mem['h13E0]=8'h46; mem['h13E1]=8'h0B; mem['h13E2]=8'h11; mem['h13E3]=8'h46;
    mem['h13E4]=8'h34; mem['h13E5]=8'h10; mem['h13E6]=8'h36; mem['h13E7]=8'h44;
    mem['h13E8]=8'hC7; mem['h13E9]=8'hA0; mem['h13EA]=8'h36; mem['h13EB]=8'h6F;
    mem['h13EC]=8'h68; mem['h13ED]=8'hF5; mem['h13EE]=8'h13; mem['h13EF]=8'hC7;
    mem['h13F0]=8'h2C; mem['h13F1]=8'hFF; mem['h13F2]=8'h04; mem['h13F3]=8'h01;
    mem['h13F4]=8'hF8; mem['h13F5]=8'h36; mem['h13F6]=8'h46; mem['h13F7]=8'hC7;
    mem['h13F8]=8'hA0; mem['h13F9]=8'h68; mem['h13FA]=8'h00; mem['h13FB]=8'h14;
    mem['h13FC]=8'h36; mem['h13FD]=8'h45; mem['h13FE]=8'hA8; mem['h13FF]=8'h97;
    mem['h1400]=8'h36; mem['h1401]=8'h6F; mem['h1402]=8'h87; mem['h1403]=8'hF8;
    mem['h1404]=8'h70; mem['h1405]=8'h1B; mem['h1406]=8'h14; mem['h1407]=8'h2B;
    mem['h1408]=8'h36; mem['h1409]=8'h88; mem['h140A]=8'h2E; mem['h140B]=8'h01;
    mem['h140C]=8'h46; mem['h140D]=8'hBF; mem['h140E]=8'h12; mem['h140F]=8'h46;
    mem['h1410]=8'h26; mem['h1411]=8'h11; mem['h1412]=8'h36; mem['h1413]=8'h6F;
    mem['h1414]=8'hD7; mem['h1415]=8'h11; mem['h1416]=8'hFA; mem['h1417]=8'h48;
    mem['h1418]=8'h08; mem['h1419]=8'h14; mem['h141A]=8'h07; mem['h141B]=8'h36;
    mem['h141C]=8'h8C; mem['h141D]=8'h2E; mem['h141E]=8'h01; mem['h141F]=8'h46;
    mem['h1420]=8'hBF; mem['h1421]=8'h12; mem['h1422]=8'h46; mem['h1423]=8'h26;
    mem['h1424]=8'h11; mem['h1425]=8'h36; mem['h1426]=8'h6F; mem['h1427]=8'hCF;
    mem['h1428]=8'h08; mem['h1429]=8'hF9; mem['h142A]=8'h48; mem['h142B]=8'h1B;
    mem['h142C]=8'h14; mem['h142D]=8'h07; mem['h142E]=8'h46; mem['h142F]=8'hCF;
    mem['h1430]=8'h12; mem['h1431]=8'h36; mem['h1432]=8'h6B; mem['h1433]=8'hC2;
    mem['h1434]=8'h24; mem['h1435]=8'h0F; mem['h1436]=8'hF8; mem['h1437]=8'h26;
    mem['h1438]=8'h68; mem['h1439]=8'h36; mem['h143A]=8'h6C; mem['h143B]=8'hDD;
    mem['h143C]=8'h0E; mem['h143D]=8'h03; mem['h143E]=8'h46; mem['h143F]=8'h0B;
    mem['h1440]=8'h11; mem['h1441]=8'h36; mem['h1442]=8'h6C; mem['h1443]=8'h0E;
    mem['h1444]=8'h03; mem['h1445]=8'h46; mem['h1446]=8'h7F; mem['h1447]=8'h12;
    mem['h1448]=8'h36; mem['h1449]=8'h6C; mem['h144A]=8'h0E; mem['h144B]=8'h03;
    mem['h144C]=8'h46; mem['h144D]=8'h7F; mem['h144E]=8'h12; mem['h144F]=8'h26;
    mem['h1450]=8'h6C; mem['h1451]=8'h36; mem['h1452]=8'h68; mem['h1453]=8'h0E;
    mem['h1454]=8'h03; mem['h1455]=8'h46; mem['h1456]=8'h57; mem['h1457]=8'h12;
    mem['h1458]=8'h36; mem['h1459]=8'h6C; mem['h145A]=8'h0E; mem['h145B]=8'h03;
    mem['h145C]=8'h46; mem['h145D]=8'h7F; mem['h145E]=8'h12; mem['h145F]=8'h36;
    mem['h1460]=8'h6A; mem['h1461]=8'hA8; mem['h1462]=8'hF8; mem['h1463]=8'h31;
    mem['h1464]=8'hF8; mem['h1465]=8'h36; mem['h1466]=8'h6B; mem['h1467]=8'hC7;
    mem['h1468]=8'h36; mem['h1469]=8'h68; mem['h146A]=8'hF8; mem['h146B]=8'h26;
    mem['h146C]=8'h6C; mem['h146D]=8'h0E; mem['h146E]=8'h03; mem['h146F]=8'h46;
    mem['h1470]=8'h57; mem['h1471]=8'h12; mem['h1472]=8'h44; mem['h1473]=8'hDF;
    mem['h1474]=8'h12; mem['h1475]=8'h2E; mem['h1476]=8'h01; mem['h1477]=8'h36;
    mem['h1478]=8'h6F; mem['h1479]=8'h3E; mem['h147A]=8'h00; mem['h147B]=8'h36;
    mem['h147C]=8'h56; mem['h147D]=8'hC7; mem['h147E]=8'hA0; mem['h147F]=8'h70;
    mem['h1480]=8'h87; mem['h1481]=8'h14; mem['h1482]=8'h06; mem['h1483]=8'hA0;
    mem['h1484]=8'h44; mem['h1485]=8'h90; mem['h1486]=8'h14; mem['h1487]=8'h36;
    mem['h1488]=8'h54; mem['h1489]=8'h0E; mem['h148A]=8'h03; mem['h148B]=8'h46;
    mem['h148C]=8'h68; mem['h148D]=8'h12; mem['h148E]=8'h06; mem['h148F]=8'hAD;
    mem['h1490]=8'h46; mem['h1491]=8'h82; mem['h1492]=8'h03; mem['h1493]=8'h36;
    mem['h1494]=8'h48; mem['h1495]=8'hC7; mem['h1496]=8'hA0; mem['h1497]=8'h68;
    mem['h1498]=8'hAB; mem['h1499]=8'h14; mem['h149A]=8'h36; mem['h149B]=8'h57;
    mem['h149C]=8'h06; mem['h149D]=8'h17; mem['h149E]=8'hCF; mem['h149F]=8'h08;
    mem['h14A0]=8'h09; mem['h14A1]=8'h70; mem['h14A2]=8'hAB; mem['h14A3]=8'h14;
    mem['h14A4]=8'h91; mem['h14A5]=8'h70; mem['h14A6]=8'hAB; mem['h14A7]=8'h14;
    mem['h14A8]=8'h44; mem['h14A9]=8'hB9; mem['h14AA]=8'h14; mem['h14AB]=8'h36;
    mem['h14AC]=8'h48; mem['h14AD]=8'h3E; mem['h14AE]=8'h00; mem['h14AF]=8'h06;
    mem['h14B0]=8'hB0; mem['h14B1]=8'h46; mem['h14B2]=8'h82; mem['h14B3]=8'h03;
    mem['h14B4]=8'h06; mem['h14B5]=8'hAE; mem['h14B6]=8'h46; mem['h14B7]=8'h82;
    mem['h14B8]=8'h03; mem['h14B9]=8'h36; mem['h14BA]=8'h57; mem['h14BB]=8'h06;
    mem['h14BC]=8'hFF; mem['h14BD]=8'h87; mem['h14BE]=8'hF8; mem['h14BF]=8'h50;
    mem['h14C0]=8'hDE; mem['h14C1]=8'h14; mem['h14C2]=8'h06; mem['h14C3]=8'h04;
    mem['h14C4]=8'h87; mem['h14C5]=8'h50; mem['h14C6]=8'hF0; mem['h14C7]=8'h14;
    mem['h14C8]=8'h36; mem['h14C9]=8'h88; mem['h14CA]=8'h2E; mem['h14CB]=8'h01;
    mem['h14CC]=8'h46; mem['h14CD]=8'hBF; mem['h14CE]=8'h12; mem['h14CF]=8'h46;
    mem['h14D0]=8'h26; mem['h14D1]=8'h11; mem['h14D2]=8'h36; mem['h14D3]=8'h6F;
    mem['h14D4]=8'hD7; mem['h14D5]=8'h11; mem['h14D6]=8'hFA; mem['h14D7]=8'h36;
    mem['h14D8]=8'h57; mem['h14D9]=8'hC7; mem['h14DA]=8'hA0; mem['h14DB]=8'h44;
    mem['h14DC]=8'hBF; mem['h14DD]=8'h14; mem['h14DE]=8'h36; mem['h14DF]=8'h8C;
    mem['h14E0]=8'h2E; mem['h14E1]=8'h01; mem['h14E2]=8'h46; mem['h14E3]=8'hBF;
    mem['h14E4]=8'h12; mem['h14E5]=8'h46; mem['h14E6]=8'h26; mem['h14E7]=8'h11;
    mem['h14E8]=8'h36; mem['h14E9]=8'h6F; mem['h14EA]=8'hCF; mem['h14EB]=8'h08;
    mem['h14EC]=8'hF9; mem['h14ED]=8'h44; mem['h14EE]=8'hD7; mem['h14EF]=8'h14;
    mem['h14F0]=8'h26; mem['h14F1]=8'h74; mem['h14F2]=8'hDD; mem['h14F3]=8'h36;
    mem['h14F4]=8'h54; mem['h14F5]=8'h0E; mem['h14F6]=8'h03; mem['h14F7]=8'h46;
    mem['h14F8]=8'h0B; mem['h14F9]=8'h11; mem['h14FA]=8'h36; mem['h14FB]=8'h77;
    mem['h14FC]=8'h3E; mem['h14FD]=8'h00; mem['h14FE]=8'h36; mem['h14FF]=8'h74;
    mem['h1500]=8'h0E; mem['h1501]=8'h03; mem['h1502]=8'h46; mem['h1503]=8'h7F;
    mem['h1504]=8'h12; mem['h1505]=8'h46; mem['h1506]=8'h93; mem['h1507]=8'h15;
    mem['h1508]=8'h36; mem['h1509]=8'h57; mem['h150A]=8'hCF; mem['h150B]=8'h08;
    mem['h150C]=8'hF9; mem['h150D]=8'h68; mem['h150E]=8'h1A; mem['h150F]=8'h15;
    mem['h1510]=8'h36; mem['h1511]=8'h77; mem['h1512]=8'h0E; mem['h1513]=8'h04;
    mem['h1514]=8'h46; mem['h1515]=8'h89; mem['h1516]=8'h12; mem['h1517]=8'h44;
    mem['h1518]=8'h08; mem['h1519]=8'h15; mem['h151A]=8'h36; mem['h151B]=8'h47;
    mem['h151C]=8'h3E; mem['h151D]=8'h07; mem['h151E]=8'h36; mem['h151F]=8'h77;
    mem['h1520]=8'hC7; mem['h1521]=8'hA0; mem['h1522]=8'h68; mem['h1523]=8'h75;
    mem['h1524]=8'h15; mem['h1525]=8'h36; mem['h1526]=8'h77; mem['h1527]=8'hC7;
    mem['h1528]=8'hA0; mem['h1529]=8'h48; mem['h152A]=8'h45; mem['h152B]=8'h15;
    mem['h152C]=8'h36; mem['h152D]=8'h48; mem['h152E]=8'hC7; mem['h152F]=8'hA0;
    mem['h1530]=8'h68; mem['h1531]=8'h44; mem['h1532]=8'h15; mem['h1533]=8'h36;
    mem['h1534]=8'h6F; mem['h1535]=8'hD7; mem['h1536]=8'h11; mem['h1537]=8'h10;
    mem['h1538]=8'h50; mem['h1539]=8'h44; mem['h153A]=8'h15; mem['h153B]=8'h36;
    mem['h153C]=8'h76; mem['h153D]=8'hC7; mem['h153E]=8'h24; mem['h153F]=8'hE0;
    mem['h1540]=8'h48; mem['h1541]=8'h44; mem['h1542]=8'h15; mem['h1543]=8'h07;
    mem['h1544]=8'hA8; mem['h1545]=8'h04; mem['h1546]=8'hB0; mem['h1547]=8'h46;
    mem['h1548]=8'h82; mem['h1549]=8'h03; mem['h154A]=8'h36; mem['h154B]=8'h48;
    mem['h154C]=8'hC7; mem['h154D]=8'hA0; mem['h154E]=8'h48; mem['h154F]=8'h5F;
    mem['h1550]=8'h15; mem['h1551]=8'h36; mem['h1552]=8'h47; mem['h1553]=8'hD7;
    mem['h1554]=8'h11; mem['h1555]=8'hFA; mem['h1556]=8'h68; mem['h1557]=8'hC0;
    mem['h1558]=8'h15; mem['h1559]=8'h46; mem['h155A]=8'h93; mem['h155B]=8'h15;
    mem['h155C]=8'h44; mem['h155D]=8'h25; mem['h155E]=8'h15; mem['h155F]=8'h36;
    mem['h1560]=8'h6F; mem['h1561]=8'hD7; mem['h1562]=8'h11; mem['h1563]=8'hFA;
    mem['h1564]=8'h48; mem['h1565]=8'h6C; mem['h1566]=8'h15; mem['h1567]=8'h06;
    mem['h1568]=8'hAE; mem['h1569]=8'h46; mem['h156A]=8'h82; mem['h156B]=8'h03;
    mem['h156C]=8'h36; mem['h156D]=8'h47; mem['h156E]=8'hD7; mem['h156F]=8'h11;
    mem['h1570]=8'hFA; mem['h1571]=8'h2B; mem['h1572]=8'h44; mem['h1573]=8'h59;
    mem['h1574]=8'h15; mem['h1575]=8'h36; mem['h1576]=8'h6F; mem['h1577]=8'hD7;
    mem['h1578]=8'h11; mem['h1579]=8'hFA; mem['h157A]=8'h36; mem['h157B]=8'h76;
    mem['h157C]=8'hC7; mem['h157D]=8'hA0; mem['h157E]=8'h48; mem['h157F]=8'h4A;
    mem['h1580]=8'h15; mem['h1581]=8'h31; mem['h1582]=8'hC7; mem['h1583]=8'hA0;
    mem['h1584]=8'h48; mem['h1585]=8'h4A; mem['h1586]=8'h15; mem['h1587]=8'h31;
    mem['h1588]=8'hC7; mem['h1589]=8'hA0; mem['h158A]=8'h48; mem['h158B]=8'h4A;
    mem['h158C]=8'h15; mem['h158D]=8'h36; mem['h158E]=8'h6F; mem['h158F]=8'hF8;
    mem['h1590]=8'h44; mem['h1591]=8'h4A; mem['h1592]=8'h15; mem['h1593]=8'h36;
    mem['h1594]=8'h77; mem['h1595]=8'h3E; mem['h1596]=8'h00; mem['h1597]=8'h36;
    mem['h1598]=8'h74; mem['h1599]=8'hDD; mem['h159A]=8'h26; mem['h159B]=8'h70;
    mem['h159C]=8'h0E; mem['h159D]=8'h04; mem['h159E]=8'h46; mem['h159F]=8'h0B;
    mem['h15A0]=8'h11; mem['h15A1]=8'h36; mem['h15A2]=8'h74; mem['h15A3]=8'h0E;
    mem['h15A4]=8'h04; mem['h15A5]=8'h46; mem['h15A6]=8'h7F; mem['h15A7]=8'h12;
    mem['h15A8]=8'h36; mem['h15A9]=8'h74; mem['h15AA]=8'h0E; mem['h15AB]=8'h04;
    mem['h15AC]=8'h46; mem['h15AD]=8'h7F; mem['h15AE]=8'h12; mem['h15AF]=8'h36;
    mem['h15B0]=8'h70; mem['h15B1]=8'h26; mem['h15B2]=8'h74; mem['h15B3]=8'h0E;
    mem['h15B4]=8'h04; mem['h15B5]=8'h46; mem['h15B6]=8'h57; mem['h15B7]=8'h12;
    mem['h15B8]=8'h36; mem['h15B9]=8'h74; mem['h15BA]=8'h0E; mem['h15BB]=8'h04;
    mem['h15BC]=8'h46; mem['h15BD]=8'h7F; mem['h15BE]=8'h12; mem['h15BF]=8'h07;
    mem['h15C0]=8'h36; mem['h15C1]=8'h6F; mem['h15C2]=8'hC7; mem['h15C3]=8'hA0;
    mem['h15C4]=8'h2B; mem['h15C5]=8'h06; mem['h15C6]=8'hC5; mem['h15C7]=8'h46;
    mem['h15C8]=8'h82; mem['h15C9]=8'h03; mem['h15CA]=8'hC7; mem['h15CB]=8'hA0;
    mem['h15CC]=8'h70; mem['h15CD]=8'hD4; mem['h15CE]=8'h15; mem['h15CF]=8'h06;
    mem['h15D0]=8'hAB; mem['h15D1]=8'h44; mem['h15D2]=8'hDB; mem['h15D3]=8'h15;
    mem['h15D4]=8'h2C; mem['h15D5]=8'hFF; mem['h15D6]=8'h04; mem['h15D7]=8'h01;
    mem['h15D8]=8'hF8; mem['h15D9]=8'h06; mem['h15DA]=8'hAD; mem['h15DB]=8'h46;
    mem['h15DC]=8'h82; mem['h15DD]=8'h03; mem['h15DE]=8'h0E; mem['h15DF]=8'h00;
    mem['h15E0]=8'hC7; mem['h15E1]=8'h14; mem['h15E2]=8'h0A; mem['h15E3]=8'h70;
    mem['h15E4]=8'hEB; mem['h15E5]=8'h15; mem['h15E6]=8'hF8; mem['h15E7]=8'h08;
    mem['h15E8]=8'h44; mem['h15E9]=8'hE1; mem['h15EA]=8'h15; mem['h15EB]=8'h06;
    mem['h15EC]=8'hB0; mem['h15ED]=8'h81; mem['h15EE]=8'h46; mem['h15EF]=8'h82;
    mem['h15F0]=8'h03; mem['h15F1]=8'hC7; mem['h15F2]=8'h04; mem['h15F3]=8'hB0;
    mem['h15F4]=8'h46; mem['h15F5]=8'h82; mem['h15F6]=8'h03; mem['h15F7]=8'h07;
    mem['h15F8]=8'hFF; mem['h15F9]=8'hFF; mem['h15FA]=8'hFF; mem['h15FB]=8'hFF;
    mem['h15FC]=8'hFF; mem['h15FD]=8'hFF; mem['h15FE]=8'hFF; mem['h15FF]=8'hFF;
    mem['h1600]=8'h00; mem['h1601]=8'hFF; mem['h1602]=8'hFF; mem['h1603]=8'hFF;
    mem['h1604]=8'hFF; mem['h1605]=8'hFF; mem['h1606]=8'hFF; mem['h1607]=8'hFF;
    mem['h1608]=8'hFF; mem['h1609]=8'hFF; mem['h160A]=8'hFF; mem['h160B]=8'hFF;
    mem['h160C]=8'hFF; mem['h160D]=8'hFF; mem['h160E]=8'hFF; mem['h160F]=8'hFF;
    mem['h1610]=8'hFF; mem['h1611]=8'hFF; mem['h1612]=8'hFF; mem['h1613]=8'hFF;
    mem['h1614]=8'hFF; mem['h1615]=8'hFF; mem['h1616]=8'hFF; mem['h1617]=8'hFF;
    mem['h1618]=8'hFF; mem['h1619]=8'hFF; mem['h161A]=8'hFF; mem['h161B]=8'hFF;
    mem['h161C]=8'hFF; mem['h161D]=8'hFF; mem['h161E]=8'hFF; mem['h161F]=8'hFF;
    mem['h1620]=8'hFF; mem['h1621]=8'hFF; mem['h1622]=8'hFF; mem['h1623]=8'hFF;
    mem['h1624]=8'hFF; mem['h1625]=8'hFF; mem['h1626]=8'hFF; mem['h1627]=8'hFF;
    mem['h1628]=8'hFF; mem['h1629]=8'hFF; mem['h162A]=8'hFF; mem['h162B]=8'hFF;
    mem['h162C]=8'hFF; mem['h162D]=8'hFF; mem['h162E]=8'hFF; mem['h162F]=8'hFF;
    mem['h1630]=8'hFF; mem['h1631]=8'hFF; mem['h1632]=8'hFF; mem['h1633]=8'hFF;
    mem['h1634]=8'hFF; mem['h1635]=8'hFF; mem['h1636]=8'hFF; mem['h1637]=8'hFF;
    mem['h1638]=8'hFF; mem['h1639]=8'hFF; mem['h163A]=8'hFF; mem['h163B]=8'hFF;
    mem['h163C]=8'hFF; mem['h163D]=8'hFF; mem['h163E]=8'hFF; mem['h163F]=8'hFF;
    mem['h1640]=8'hFF; mem['h1641]=8'hFF; mem['h1642]=8'hFF; mem['h1643]=8'hFF;
    mem['h1644]=8'hFF; mem['h1645]=8'hFF; mem['h1646]=8'hFF; mem['h1647]=8'hFF;
    mem['h1648]=8'hFF; mem['h1649]=8'hFF; mem['h164A]=8'hFF; mem['h164B]=8'hFF;
    mem['h164C]=8'hFF; mem['h164D]=8'hFF; mem['h164E]=8'hFF; mem['h164F]=8'hFF;
    mem['h1650]=8'h00; mem['h1651]=8'h00; mem['h1652]=8'h00; mem['h1653]=8'h00;
    mem['h1654]=8'h00; mem['h1655]=8'h00; mem['h1656]=8'h00; mem['h1657]=8'h00;
    mem['h1658]=8'h00; mem['h1659]=8'h00; mem['h165A]=8'h00; mem['h165B]=8'h00;
    mem['h165C]=8'h00; mem['h165D]=8'h00; mem['h165E]=8'h00; mem['h165F]=8'h00;
    mem['h1660]=8'h00; mem['h1661]=8'h00; mem['h1662]=8'h00; mem['h1663]=8'h00;
    mem['h1664]=8'h00; mem['h1665]=8'h00; mem['h1666]=8'h00; mem['h1667]=8'h00;
    mem['h1668]=8'h00; mem['h1669]=8'h00; mem['h166A]=8'h00; mem['h166B]=8'h00;
    mem['h166C]=8'h00; mem['h166D]=8'h00; mem['h166E]=8'h00; mem['h166F]=8'h00;
    mem['h1670]=8'h00; mem['h1671]=8'h00; mem['h1672]=8'h00; mem['h1673]=8'h00;
    mem['h1674]=8'h00; mem['h1675]=8'h00; mem['h1676]=8'h00; mem['h1677]=8'h00;
    mem['h1678]=8'h00; mem['h1679]=8'h00; mem['h167A]=8'h00; mem['h167B]=8'h00;
    mem['h167C]=8'h00; mem['h167D]=8'h00; mem['h167E]=8'h00; mem['h167F]=8'h00;
    mem['h1680]=8'h00; mem['h1681]=8'h00; mem['h1682]=8'h00; mem['h1683]=8'h00;
    mem['h1684]=8'h00; mem['h1685]=8'h00; mem['h1686]=8'h00; mem['h1687]=8'h00;
    mem['h1688]=8'h00; mem['h1689]=8'hFF; mem['h168A]=8'hFF; mem['h168B]=8'hFF;
    mem['h168C]=8'hFF; mem['h168D]=8'hFF; mem['h168E]=8'hFF; mem['h168F]=8'hFF;
    mem['h1690]=8'hFF; mem['h1691]=8'hFF; mem['h1692]=8'hFF; mem['h1693]=8'hFF;
    mem['h1694]=8'hFF; mem['h1695]=8'hFF; mem['h1696]=8'hFF; mem['h1697]=8'hFF;
    mem['h1698]=8'h00; mem['h1699]=8'hFF; mem['h169A]=8'hFF; mem['h169B]=8'hFF;
    mem['h169C]=8'hFF; mem['h169D]=8'hFF; mem['h169E]=8'hFF; mem['h169F]=8'hFF;
    mem['h16A0]=8'h00; mem['h16A1]=8'h03; mem['h16A2]=8'h03; mem['h16A3]=8'h04;
    mem['h16A4]=8'h04; mem['h16A5]=8'h05; mem['h16A6]=8'h06; mem['h16A7]=8'h01;
    mem['h16A8]=8'h02; mem['h16A9]=8'h02; mem['h16AA]=8'h02; mem['h16AB]=8'h02;
    mem['h16AC]=8'h02; mem['h16AD]=8'h02; mem['h16AE]=8'h02; mem['h16AF]=8'h00;
    mem['h16B0]=8'h03; mem['h16B1]=8'h03; mem['h16B2]=8'h04; mem['h16B3]=8'h04;
    mem['h16B4]=8'h05; mem['h16B5]=8'h01; mem['h16B6]=8'h01; mem['h16B7]=8'h02;
    mem['h16B8]=8'h02; mem['h16B9]=8'h02; mem['h16BA]=8'h02; mem['h16BB]=8'h02;
    mem['h16BC]=8'h02; mem['h16BD]=8'h02; mem['h16BE]=8'h00; mem['h16BF]=8'h00;
    mem['h16C0]=8'h03; mem['h16C1]=8'hC9; mem['h16C2]=8'hCE; mem['h16C3]=8'hD4;
    mem['h16C4]=8'h03; mem['h16C5]=8'hD3; mem['h16C6]=8'hC7; mem['h16C7]=8'hCE;
    mem['h16C8]=8'h03; mem['h16C9]=8'hC1; mem['h16CA]=8'hC2; mem['h16CB]=8'hD3;
    mem['h16CC]=8'h03; mem['h16CD]=8'hD3; mem['h16CE]=8'hD1; mem['h16CF]=8'hD2;
    mem['h16D0]=8'h03; mem['h16D1]=8'hD4; mem['h16D2]=8'hC1; mem['h16D3]=8'hC2;
    mem['h16D4]=8'h03; mem['h16D5]=8'hD2; mem['h16D6]=8'hCE; mem['h16D7]=8'hC4;
    mem['h16D8]=8'h03; mem['h16D9]=8'hC3; mem['h16DA]=8'hC8; mem['h16DB]=8'hD2;
    mem['h16DC]=8'h03; mem['h16DD]=8'hD5; mem['h16DE]=8'hC4; mem['h16DF]=8'hC6;
    mem['h16E0]=8'h00; mem['h16E1]=8'h00; mem['h16E2]=8'h00; mem['h16E3]=8'h00;
    mem['h16E4]=8'h00; mem['h16E5]=8'h00; mem['h16E6]=8'h00; mem['h16E7]=8'h00;
    mem['h16E8]=8'h00; mem['h16E9]=8'h00; mem['h16EA]=8'h00; mem['h16EB]=8'h00;
    mem['h16EC]=8'h00; mem['h16ED]=8'h00; mem['h16EE]=8'h00; mem['h16EF]=8'h00;
    mem['h16F0]=8'h1B; mem['h16F1]=8'h00; mem['h16F2]=8'h00; mem['h16F3]=8'h00;
    mem['h16F4]=8'h00; mem['h16F5]=8'h00; mem['h16F6]=8'h00; mem['h16F7]=8'h00;
    mem['h16F8]=8'h00; mem['h16F9]=8'hFF; mem['h16FA]=8'hFF; mem['h16FB]=8'hFF;
    mem['h16FC]=8'hFF; mem['h16FD]=8'hFF; mem['h16FE]=8'hFF; mem['h16FF]=8'hFF;
    mem['h1700]=8'h03; mem['h1701]=8'hD2; mem['h1702]=8'hC5; mem['h1703]=8'hCD;
    mem['h1704]=8'h02; mem['h1705]=8'hC9; mem['h1706]=8'hC6; mem['h1707]=8'h03;
    mem['h1708]=8'hCC; mem['h1709]=8'hC5; mem['h170A]=8'hD4; mem['h170B]=8'h04;
    mem['h170C]=8'hC7; mem['h170D]=8'hCF; mem['h170E]=8'hD4; mem['h170F]=8'hCF;
    mem['h1710]=8'h05; mem['h1711]=8'hD0; mem['h1712]=8'hD2; mem['h1713]=8'hC9;
    mem['h1714]=8'hCE; mem['h1715]=8'hD4; mem['h1716]=8'h05; mem['h1717]=8'hC9;
    mem['h1718]=8'hCE; mem['h1719]=8'hD0; mem['h171A]=8'hD5; mem['h171B]=8'hD4;
    mem['h171C]=8'h03; mem['h171D]=8'hC6; mem['h171E]=8'hCF; mem['h171F]=8'hD2;
    mem['h1720]=8'h04; mem['h1721]=8'hCE; mem['h1722]=8'hC5; mem['h1723]=8'hD8;
    mem['h1724]=8'hD4; mem['h1725]=8'h05; mem['h1726]=8'hC7; mem['h1727]=8'hCF;
    mem['h1728]=8'hD3; mem['h1729]=8'hD5; mem['h172A]=8'hC2; mem['h172B]=8'h06;
    mem['h172C]=8'hD2; mem['h172D]=8'hC5; mem['h172E]=8'hD4; mem['h172F]=8'hD5;
    mem['h1730]=8'hD2; mem['h1731]=8'hCE; mem['h1732]=8'h03; mem['h1733]=8'hC4;
    mem['h1734]=8'hC9; mem['h1735]=8'hCD; mem['h1736]=8'h03; mem['h1737]=8'hC5;
    mem['h1738]=8'hCE; mem['h1739]=8'hC4; mem['h173A]=8'h00; mem['h173B]=8'h00;
    mem['h173C]=8'hFF; mem['h173D]=8'h00; mem['h173E]=8'h00; mem['h173F]=8'h00;
    mem['h1740]=8'h00; mem['h1741]=8'h00; mem['h1742]=8'h00; mem['h1743]=8'h00;
    mem['h1744]=8'h00; mem['h1745]=8'h00; mem['h1746]=8'h00; mem['h1747]=8'h00;
    mem['h1748]=8'h00; mem['h1749]=8'h00; mem['h174A]=8'h00; mem['h174B]=8'h00;
    mem['h174C]=8'h00; mem['h174D]=8'h00; mem['h174E]=8'h00; mem['h174F]=8'h00;
    mem['h1750]=8'h00; mem['h1751]=8'h00; mem['h1752]=8'h00; mem['h1753]=8'h00;
    mem['h1754]=8'h00; mem['h1755]=8'h00; mem['h1756]=8'h00; mem['h1757]=8'h00;
    mem['h1758]=8'h00; mem['h1759]=8'h00; mem['h175A]=8'h00; mem['h175B]=8'h00;
    mem['h175C]=8'h00; mem['h175D]=8'h00; mem['h175E]=8'h00; mem['h175F]=8'h00;
    mem['h1760]=8'h00; mem['h1761]=8'h00; mem['h1762]=8'h00; mem['h1763]=8'h00;
    mem['h1764]=8'h00; mem['h1765]=8'h00; mem['h1766]=8'h00; mem['h1767]=8'h00;
    mem['h1768]=8'h00; mem['h1769]=8'h00; mem['h176A]=8'h00; mem['h176B]=8'h00;
    mem['h176C]=8'h00; mem['h176D]=8'h00; mem['h176E]=8'h00; mem['h176F]=8'h00;
    mem['h1770]=8'h00; mem['h1771]=8'h00; mem['h1772]=8'h00; mem['h1773]=8'h00;
    mem['h1774]=8'h00; mem['h1775]=8'h00; mem['h1776]=8'h00; mem['h1777]=8'h00;
    mem['h1778]=8'h00; mem['h1779]=8'h00; mem['h177A]=8'h00; mem['h177B]=8'h00;
    mem['h177C]=8'h00; mem['h177D]=8'h00; mem['h177E]=8'h00; mem['h177F]=8'h00;
    mem['h1780]=8'h00; mem['h1781]=8'h00; mem['h1782]=8'h00; mem['h1783]=8'h00;
    mem['h1784]=8'h00; mem['h1785]=8'hFF; mem['h1786]=8'hFF; mem['h1787]=8'hFF;
    mem['h1788]=8'h00; mem['h1789]=8'hFF; mem['h178A]=8'hFF; mem['h178B]=8'hFF;
    mem['h178C]=8'hFF; mem['h178D]=8'hFF; mem['h178E]=8'hFF; mem['h178F]=8'hFF;
    mem['h1790]=8'hFF; mem['h1791]=8'hFF; mem['h1792]=8'hFF; mem['h1793]=8'hFF;
    mem['h1794]=8'hFF; mem['h1795]=8'hFF; mem['h1796]=8'hFF; mem['h1797]=8'hFF;
    mem['h1798]=8'hFF; mem['h1799]=8'hFF; mem['h179A]=8'hFF; mem['h179B]=8'hFF;
    mem['h179C]=8'hFF; mem['h179D]=8'hFF; mem['h179E]=8'hFF; mem['h179F]=8'hFF;
    mem['h17A0]=8'hFF; mem['h17A1]=8'hFF; mem['h17A2]=8'hFF; mem['h17A3]=8'hFF;
    mem['h17A4]=8'hFF; mem['h17A5]=8'hFF; mem['h17A6]=8'hFF; mem['h17A7]=8'hFF;
    mem['h17A8]=8'hFF; mem['h17A9]=8'hFF; mem['h17AA]=8'hFF; mem['h17AB]=8'hFF;
    mem['h17AC]=8'hFF; mem['h17AD]=8'hFF; mem['h17AE]=8'hFF; mem['h17AF]=8'hFF;
    mem['h17B0]=8'hFF; mem['h17B1]=8'hFF; mem['h17B2]=8'hFF; mem['h17B3]=8'hFF;
    mem['h17B4]=8'hFF; mem['h17B5]=8'hFF; mem['h17B6]=8'hFF; mem['h17B7]=8'hFF;
    mem['h17B8]=8'hFF; mem['h17B9]=8'hFF; mem['h17BA]=8'hFF; mem['h17BB]=8'hFF;
    mem['h17BC]=8'hFF; mem['h17BD]=8'hFF; mem['h17BE]=8'hFF; mem['h17BF]=8'hFF;
    mem['h17C0]=8'hFF; mem['h17C1]=8'hFF; mem['h17C2]=8'hFF; mem['h17C3]=8'hFF;
    mem['h17C4]=8'hFF; mem['h17C5]=8'hFF; mem['h17C6]=8'hFF; mem['h17C7]=8'hFF;
    mem['h17C8]=8'hFF; mem['h17C9]=8'hFF; mem['h17CA]=8'hFF; mem['h17CB]=8'hFF;
    mem['h17CC]=8'hFF; mem['h17CD]=8'hFF; mem['h17CE]=8'hFF; mem['h17CF]=8'hFF;
    mem['h17D0]=8'hFF; mem['h17D1]=8'hFF; mem['h17D2]=8'hFF; mem['h17D3]=8'hFF;
    mem['h17D4]=8'hFF; mem['h17D5]=8'hFF; mem['h17D6]=8'hFF; mem['h17D7]=8'hFF;
    mem['h17D8]=8'hFF; mem['h17D9]=8'hFF; mem['h17DA]=8'hFF; mem['h17DB]=8'hFF;
    mem['h17DC]=8'hFF; mem['h17DD]=8'hFF; mem['h17DE]=8'hFF; mem['h17DF]=8'hFF;
    mem['h17E0]=8'hFF; mem['h17E1]=8'hFF; mem['h17E2]=8'hFF; mem['h17E3]=8'hFF;
    mem['h17E4]=8'hFF; mem['h17E5]=8'hFF; mem['h17E6]=8'hFF; mem['h17E7]=8'hFF;
    mem['h17E8]=8'hFF; mem['h17E9]=8'hFF; mem['h17EA]=8'hFF; mem['h17EB]=8'hFF;
    mem['h17EC]=8'hFF; mem['h17ED]=8'hFF; mem['h17EE]=8'hFF; mem['h17EF]=8'hFF;
    mem['h17F0]=8'hFF; mem['h17F1]=8'hFF; mem['h17F2]=8'hFF; mem['h17F3]=8'hFF;
    mem['h17F4]=8'hFF; mem['h17F5]=8'hFF; mem['h17F6]=8'hFF; mem['h17F7]=8'hFF;
    mem['h17F8]=8'hFF; mem['h17F9]=8'hFF; mem['h17FA]=8'hFF; mem['h17FB]=8'hFF;
    mem['h17FC]=8'hFF; mem['h17FD]=8'hFF; mem['h17FE]=8'hFF; mem['h17FF]=8'hFF;
    mem['h1800]=8'h36; mem['h1801]=8'h53; mem['h1802]=8'h3E; mem['h1803]=8'h00;
    mem['h1804]=8'h36; mem['h1805]=8'h5B; mem['h1806]=8'h3E; mem['h1807]=8'h00;
    mem['h1808]=8'h07; mem['h1809]=8'hFF; mem['h180A]=8'hFF; mem['h180B]=8'h36;
    mem['h180C]=8'h64; mem['h180D]=8'h2E; mem['h180E]=8'h16; mem['h180F]=8'h3E;
    mem['h1810]=8'h00; mem['h1811]=8'h36; mem['h1812]=8'h82; mem['h1813]=8'hCF;
    mem['h1814]=8'h08; mem['h1815]=8'h36; mem['h1816]=8'h81; mem['h1817]=8'hF9;
    mem['h1818]=8'h36; mem['h1819]=8'h81; mem['h181A]=8'h46; mem['h181B]=8'hA0;
    mem['h181C]=8'h02; mem['h181D]=8'h68; mem['h181E]=8'h25; mem['h181F]=8'h18;
    mem['h1820]=8'h36; mem['h1821]=8'h64; mem['h1822]=8'h46; mem['h1823]=8'hCC;
    mem['h1824]=8'h02; mem['h1825]=8'h36; mem['h1826]=8'h81; mem['h1827]=8'h46;
    mem['h1828]=8'h03; mem['h1829]=8'h03; mem['h182A]=8'h48; mem['h182B]=8'h18;
    mem['h182C]=8'h18; mem['h182D]=8'h36; mem['h182E]=8'h64; mem['h182F]=8'hC7;
    mem['h1830]=8'h3C; mem['h1831]=8'h01; mem['h1832]=8'h48; mem['h1833]=8'h39;
    mem['h1834]=8'h18; mem['h1835]=8'h36; mem['h1836]=8'h66; mem['h1837]=8'h3E;
    mem['h1838]=8'h00; mem['h1839]=8'h36; mem['h183A]=8'h85; mem['h183B]=8'h2E;
    mem['h183C]=8'h17; mem['h183D]=8'hC7; mem['h183E]=8'h02; mem['h183F]=8'h02;
    mem['h1840]=8'h04; mem['h1841]=8'h5E; mem['h1842]=8'h2E; mem['h1843]=8'h17;
    mem['h1844]=8'hF0; mem['h1845]=8'h1E; mem['h1846]=8'h16; mem['h1847]=8'h26;
    mem['h1848]=8'h65; mem['h1849]=8'h0E; mem['h184A]=8'h02; mem['h184B]=8'h46;
    mem['h184C]=8'hF8; mem['h184D]=8'h02; mem['h184E]=8'h68; mem['h184F]=8'h58;
    mem['h1850]=8'h18; mem['h1851]=8'h06; mem['h1852]=8'hC6; mem['h1853]=8'h16;
    mem['h1854]=8'hCE; mem['h1855]=8'h44; mem['h1856]=8'h96; mem['h1857]=8'h02;
    mem['h1858]=8'h36; mem['h1859]=8'hF0; mem['h185A]=8'h2E; mem['h185B]=8'h16;
    mem['h185C]=8'hDF; mem['h185D]=8'h30; mem['h185E]=8'hE7; mem['h185F]=8'h30;
    mem['h1860]=8'hFB; mem['h1861]=8'h30; mem['h1862]=8'hFC; mem['h1863]=8'h36;
    mem['h1864]=8'h85; mem['h1865]=8'h2E; mem['h1866]=8'h17; mem['h1867]=8'hC7;
    mem['h1868]=8'h02; mem['h1869]=8'h02; mem['h186A]=8'h04; mem['h186B]=8'h5C;
    mem['h186C]=8'hF0; mem['h186D]=8'hDF; mem['h186E]=8'h30; mem['h186F]=8'hE7;
    mem['h1870]=8'h36; mem['h1871]=8'hF0; mem['h1872]=8'h2E; mem['h1873]=8'h16;
    mem['h1874]=8'hFB; mem['h1875]=8'h30; mem['h1876]=8'hFC; mem['h1877]=8'hEB;
    mem['h1878]=8'hF4; mem['h1879]=8'h1E; mem['h187A]=8'h16; mem['h187B]=8'h26;
    mem['h187C]=8'h00; mem['h187D]=8'h46; mem['h187E]=8'h26; mem['h187F]=8'h0A;
    mem['h1880]=8'h36; mem['h1881]=8'hD5; mem['h1882]=8'h2E; mem['h1883]=8'h01;
    mem['h1884]=8'h46; mem['h1885]=8'h0A; mem['h1886]=8'h0B; mem['h1887]=8'hC4;
    mem['h1888]=8'hA0; mem['h1889]=8'h68; mem['h188A]=8'h51; mem['h188B]=8'h18;
    mem['h188C]=8'h04; mem['h188D]=8'h02; mem['h188E]=8'h36; mem['h188F]=8'hBE;
    mem['h1890]=8'h2E; mem['h1891]=8'h16; mem['h1892]=8'hF8; mem['h1893]=8'h36;
    mem['h1894]=8'hD8; mem['h1895]=8'h2E; mem['h1896]=8'h01; mem['h1897]=8'h46;
    mem['h1898]=8'h0A; mem['h1899]=8'h0B; mem['h189A]=8'hC4; mem['h189B]=8'hA0;
    mem['h189C]=8'h48; mem['h189D]=8'hC0; mem['h189E]=8'h18; mem['h189F]=8'h36;
    mem['h18A0]=8'h04; mem['h18A1]=8'h2E; mem['h18A2]=8'h01; mem['h18A3]=8'h46;
    mem['h18A4]=8'hA4; mem['h18A5]=8'h12; mem['h18A6]=8'h36; mem['h18A7]=8'hC4;
    mem['h18A8]=8'h46; mem['h18A9]=8'hAD; mem['h18AA]=8'h12; mem['h18AB]=8'h36;
    mem['h18AC]=8'h00; mem['h18AD]=8'h2E; mem['h18AE]=8'h16; mem['h18AF]=8'hCF;
    mem['h18B0]=8'h36; mem['h18B1]=8'hBF; mem['h18B2]=8'hF9; mem['h18B3]=8'h46;
    mem['h18B4]=8'h94; mem['h18B5]=8'h03; mem['h18B6]=8'h36; mem['h18B7]=8'hC8;
    mem['h18B8]=8'h2E; mem['h18B9]=8'h01; mem['h18BA]=8'h46; mem['h18BB]=8'hAD;
    mem['h18BC]=8'h12; mem['h18BD]=8'h44; mem['h18BE]=8'hE9; mem['h18BF]=8'h18;
    mem['h18C0]=8'h21; mem['h18C1]=8'h36; mem['h18C2]=8'hBF; mem['h18C3]=8'h2E;
    mem['h18C4]=8'h16; mem['h18C5]=8'hFC; mem['h18C6]=8'h46; mem['h18C7]=8'h94;
    mem['h18C8]=8'h03; mem['h18C9]=8'h36; mem['h18CA]=8'hC8; mem['h18CB]=8'h2E;
    mem['h18CC]=8'h01; mem['h18CD]=8'h46; mem['h18CE]=8'hAD; mem['h18CF]=8'h12;
    mem['h18D0]=8'h36; mem['h18D1]=8'hBF; mem['h18D2]=8'h2E; mem['h18D3]=8'h16;
    mem['h18D4]=8'hC7; mem['h18D5]=8'h04; mem['h18D6]=8'h05; mem['h18D7]=8'h31;
    mem['h18D8]=8'hF8; mem['h18D9]=8'h36; mem['h18DA]=8'h00; mem['h18DB]=8'hCF;
    mem['h18DC]=8'h36; mem['h18DD]=8'hBF; mem['h18DE]=8'hF9; mem['h18DF]=8'h46;
    mem['h18E0]=8'h94; mem['h18E1]=8'h03; mem['h18E2]=8'h36; mem['h18E3]=8'hC4;
    mem['h18E4]=8'h2E; mem['h18E5]=8'h01; mem['h18E6]=8'h46; mem['h18E7]=8'hAD;
    mem['h18E8]=8'h12; mem['h18E9]=8'h36; mem['h18EA]=8'h64; mem['h18EB]=8'h2E;
    mem['h18EC]=8'h16; mem['h18ED]=8'h3E; mem['h18EE]=8'h00; mem['h18EF]=8'h36;
    mem['h18F0]=8'h1C; mem['h18F1]=8'h2E; mem['h18F2]=8'h17; mem['h18F3]=8'h46;
    mem['h18F4]=8'h0A; mem['h18F5]=8'h0B; mem['h18F6]=8'hC4; mem['h18F7]=8'hA0;
    mem['h18F8]=8'h36; mem['h18F9]=8'h82; mem['h18FA]=8'h2E; mem['h18FB]=8'h16;
    mem['h18FC]=8'hF8; mem['h18FD]=8'h68; mem['h18FE]=8'h51; mem['h18FF]=8'h18;
    mem['h1900]=8'h04; mem['h1901]=8'h03; mem['h1902]=8'h36; mem['h1903]=8'h83;
    mem['h1904]=8'hF8; mem['h1905]=8'h36; mem['h1906]=8'h83; mem['h1907]=8'h46;
    mem['h1908]=8'hA0; mem['h1909]=8'h02; mem['h190A]=8'h68; mem['h190B]=8'h17;
    mem['h190C]=8'h19; mem['h190D]=8'h3C; mem['h190E]=8'hBD; mem['h190F]=8'h68;
    mem['h1910]=8'h22; mem['h1911]=8'h19; mem['h1912]=8'h36; mem['h1913]=8'h64;
    mem['h1914]=8'h46; mem['h1915]=8'hCC; mem['h1916]=8'h02; mem['h1917]=8'h36;
    mem['h1918]=8'h83; mem['h1919]=8'h46; mem['h191A]=8'h03; mem['h191B]=8'h03;
    mem['h191C]=8'h48; mem['h191D]=8'h05; mem['h191E]=8'h19; mem['h191F]=8'h44;
    mem['h1920]=8'h51; mem['h1921]=8'h18; mem['h1922]=8'h36; mem['h1923]=8'h82;
    mem['h1924]=8'h2E; mem['h1925]=8'h16; mem['h1926]=8'hC7; mem['h1927]=8'h04;
    mem['h1928]=8'h03; mem['h1929]=8'h36; mem['h192A]=8'hBE; mem['h192B]=8'hF8;
    mem['h192C]=8'h36; mem['h192D]=8'h83; mem['h192E]=8'hCF; mem['h192F]=8'h09;
    mem['h1930]=8'h36; mem['h1931]=8'hBF; mem['h1932]=8'hF9; mem['h1933]=8'h46;
    mem['h1934]=8'h94; mem['h1935]=8'h03; mem['h1936]=8'h36; mem['h1937]=8'hC4;
    mem['h1938]=8'h2E; mem['h1939]=8'h01; mem['h193A]=8'h46; mem['h193B]=8'hBF;
    mem['h193C]=8'h12; mem['h193D]=8'h46; mem['h193E]=8'h89; mem['h193F]=8'h10;
    mem['h1940]=8'h36; mem['h1941]=8'hCC; mem['h1942]=8'h2E; mem['h1943]=8'h01;
    mem['h1944]=8'h46; mem['h1945]=8'hAD; mem['h1946]=8'h12; mem['h1947]=8'h36;
    mem['h1948]=8'hC8; mem['h1949]=8'h46; mem['h194A]=8'hBF; mem['h194B]=8'h12;
    mem['h194C]=8'h46; mem['h194D]=8'h1A; mem['h194E]=8'h11; mem['h194F]=8'h36;
    mem['h1950]=8'hC6; mem['h1951]=8'hC7; mem['h1952]=8'hA0; mem['h1953]=8'h36;
    mem['h1954]=8'h56; mem['h1955]=8'hC7; mem['h1956]=8'h68; mem['h1957]=8'h51;
    mem['h1958]=8'h18; mem['h1959]=8'h70; mem['h195A]=8'h78; mem['h195B]=8'h19;
    mem['h195C]=8'hA0; mem['h195D]=8'h70; mem['h195E]=8'h7F; mem['h195F]=8'h19;
    mem['h1960]=8'h68; mem['h1961]=8'h7F; mem['h1962]=8'h19; mem['h1963]=8'h36;
    mem['h1964]=8'hF3; mem['h1965]=8'h2E; mem['h1966]=8'h16; mem['h1967]=8'hE7;
    mem['h1968]=8'h31; mem['h1969]=8'hDF; mem['h196A]=8'h31; mem['h196B]=8'hFC;
    mem['h196C]=8'h31; mem['h196D]=8'hFB; mem['h196E]=8'h36; mem['h196F]=8'h85;
    mem['h1970]=8'h2E; mem['h1971]=8'h17; mem['h1972]=8'hCF; mem['h1973]=8'h09;
    mem['h1974]=8'hF9; mem['h1975]=8'h44; mem['h1976]=8'h4E; mem['h1977]=8'h0B;
    mem['h1978]=8'hA0; mem['h1979]=8'h50; mem['h197A]=8'h7F; mem['h197B]=8'h19;
    mem['h197C]=8'h44; mem['h197D]=8'h63; mem['h197E]=8'h19; mem['h197F]=8'h36;
    mem['h1980]=8'hCC; mem['h1981]=8'h2E; mem['h1982]=8'h01; mem['h1983]=8'h46;
    mem['h1984]=8'hA4; mem['h1985]=8'h12; mem['h1986]=8'h46; mem['h1987]=8'hAA;
    mem['h1988]=8'h08; mem['h1989]=8'h46; mem['h198A]=8'h2D; mem['h198B]=8'h08;
    mem['h198C]=8'h44; mem['h198D]=8'h4E; mem['h198E]=8'h0B; mem['h198F]=8'h06;
    mem['h1990]=8'h8D; mem['h1991]=8'h46; mem['h1992]=8'h82; mem['h1993]=8'h03;
    mem['h1994]=8'h46; mem['h1995]=8'h82; mem['h1996]=8'h03; mem['h1997]=8'h36;
    mem['h1998]=8'h23; mem['h1999]=8'h2E; mem['h199A]=8'h01; mem['h199B]=8'h3E;
    mem['h199C]=8'h01; mem['h199D]=8'h36; mem['h199E]=8'h54; mem['h199F]=8'hC7;
    mem['h19A0]=8'hA0; mem['h19A1]=8'h33; mem['h19A2]=8'h2B; mem['h19A3]=8'h44;
    mem['h19A4]=8'h12; mem['h19A5]=8'h08; mem['h19A6]=8'h36; mem['h19A7]=8'h85;
    mem['h19A8]=8'h2E; mem['h19A9]=8'h17; mem['h19AA]=8'hC7; mem['h19AB]=8'h02;
    mem['h19AC]=8'h02; mem['h19AD]=8'h04; mem['h19AE]=8'h5E; mem['h19AF]=8'hE0;
    mem['h19B0]=8'hDD; mem['h19B1]=8'h36; mem['h19B2]=8'h65; mem['h19B3]=8'h2E;
    mem['h19B4]=8'h16; mem['h19B5]=8'h0E; mem['h19B6]=8'h02; mem['h19B7]=8'h46;
    mem['h19B8]=8'h0B; mem['h19B9]=8'h11; mem['h19BA]=8'h46; mem['h19BB]=8'h2D;
    mem['h19BC]=8'h08; mem['h19BD]=8'h44; mem['h19BE]=8'h4E; mem['h19BF]=8'h0B;
    mem['h19C0]=8'h36; mem['h19C1]=8'h7E; mem['h19C2]=8'h3E; mem['h19C3]=8'h00;
    mem['h19C4]=8'h46; mem['h19C5]=8'hD4; mem['h19C6]=8'h04; mem['h19C7]=8'h36;
    mem['h19C8]=8'h97; mem['h19C9]=8'h2E; mem['h19CA]=8'h01; mem['h19CB]=8'hC7;
    mem['h19CC]=8'h3C; mem['h19CD]=8'h98; mem['h19CE]=8'h2B; mem['h19CF]=8'h44;
    mem['h19D0]=8'h6A; mem['h19D1]=8'h09; mem['h19D2]=8'hFF; mem['h19D3]=8'hFF;
    mem['h19D4]=8'hFF; mem['h19D5]=8'hFF; mem['h19D6]=8'hFF; mem['h19D7]=8'hFF;
    mem['h19D8]=8'hFF; mem['h19D9]=8'hFF; mem['h19DA]=8'hFF; mem['h19DB]=8'hFF;
    mem['h19DC]=8'hFF; mem['h19DD]=8'hFF; mem['h19DE]=8'hFF; mem['h19DF]=8'hFF;
    mem['h19E0]=8'hFF; mem['h19E1]=8'hFF; mem['h19E2]=8'hFF; mem['h19E3]=8'hFF;
    mem['h19E4]=8'hFF; mem['h19E5]=8'hFF; mem['h19E6]=8'hFF; mem['h19E7]=8'hFF;
    mem['h19E8]=8'hFF; mem['h19E9]=8'hFF; mem['h19EA]=8'hFF; mem['h19EB]=8'hFF;
    mem['h19EC]=8'hFF; mem['h19ED]=8'hFF; mem['h19EE]=8'hFF; mem['h19EF]=8'hFF;
    mem['h19F0]=8'hFF; mem['h19F1]=8'hFF; mem['h19F2]=8'hFF; mem['h19F3]=8'hFF;
    mem['h19F4]=8'hFF; mem['h19F5]=8'hFF; mem['h19F6]=8'hFF; mem['h19F7]=8'hFF;
    mem['h19F8]=8'hFF; mem['h19F9]=8'hFF; mem['h19FA]=8'hFF; mem['h19FB]=8'hFF;
    mem['h19FC]=8'hFF; mem['h19FD]=8'hFF; mem['h19FE]=8'hFF; mem['h19FF]=8'hFF;
    mem['h1A00]=8'h36; mem['h1A01]=8'h0C; mem['h1A02]=8'h2E; mem['h1A03]=8'h01;
    mem['h1A04]=8'h46; mem['h1A05]=8'hAD; mem['h1A06]=8'h12; mem['h1A07]=8'h36;
    mem['h1A08]=8'h56; mem['h1A09]=8'hC7; mem['h1A0A]=8'hA0; mem['h1A0B]=8'h70;
    mem['h1A0C]=8'h8F; mem['h1A0D]=8'h1A; mem['h1A0E]=8'h68; mem['h1A0F]=8'hA7;
    mem['h1A10]=8'h06; mem['h1A11]=8'h36; mem['h1A12]=8'h0F; mem['h1A13]=8'hC7;
    mem['h1A14]=8'hA0; mem['h1A15]=8'h70; mem['h1A16]=8'h21; mem['h1A17]=8'h1A;
    mem['h1A18]=8'h1A; mem['h1A19]=8'hC8; mem['h1A1A]=8'h06; mem['h1A1B]=8'h00;
    mem['h1A1C]=8'h12; mem['h1A1D]=8'hF8; mem['h1A1E]=8'h44; mem['h1A1F]=8'h32;
    mem['h1A20]=8'h1A; mem['h1A21]=8'hC8; mem['h1A22]=8'hA8; mem['h1A23]=8'h91;
    mem['h1A24]=8'hA0; mem['h1A25]=8'h1A; mem['h1A26]=8'hC8; mem['h1A27]=8'h06;
    mem['h1A28]=8'h00; mem['h1A29]=8'h88; mem['h1A2A]=8'hF8; mem['h1A2B]=8'h68;
    mem['h1A2C]=8'h2F; mem['h1A2D]=8'h1A; mem['h1A2E]=8'h08; mem['h1A2F]=8'hA8;
    mem['h1A30]=8'h91; mem['h1A31]=8'hC8; mem['h1A32]=8'h36; mem['h1A33]=8'h0B;
    mem['h1A34]=8'hF9; mem['h1A35]=8'h36; mem['h1A36]=8'h04; mem['h1A37]=8'h26;
    mem['h1A38]=8'h1C; mem['h1A39]=8'hDD; mem['h1A3A]=8'h0E; mem['h1A3B]=8'h04;
    mem['h1A3C]=8'h46; mem['h1A3D]=8'h0B; mem['h1A3E]=8'h11; mem['h1A3F]=8'h46;
    mem['h1A40]=8'hA7; mem['h1A41]=8'h06; mem['h1A42]=8'h36; mem['h1A43]=8'h24;
    mem['h1A44]=8'h46; mem['h1A45]=8'hAD; mem['h1A46]=8'h12; mem['h1A47]=8'h36;
    mem['h1A48]=8'h1C; mem['h1A49]=8'h46; mem['h1A4A]=8'hA4; mem['h1A4B]=8'h12;
    mem['h1A4C]=8'h36; mem['h1A4D]=8'h0C; mem['h1A4E]=8'h46; mem['h1A4F]=8'hB6;
    mem['h1A50]=8'h12; mem['h1A51]=8'h46; mem['h1A52]=8'hD2; mem['h1A53]=8'h11;
    mem['h1A54]=8'h36; mem['h1A55]=8'h1C; mem['h1A56]=8'h46; mem['h1A57]=8'hB6;
    mem['h1A58]=8'h12; mem['h1A59]=8'h46; mem['h1A5A]=8'h89; mem['h1A5B]=8'h10;
    mem['h1A5C]=8'h36; mem['h1A5D]=8'h57; mem['h1A5E]=8'hCF; mem['h1A5F]=8'h09;
    mem['h1A60]=8'hF9; mem['h1A61]=8'h36; mem['h1A62]=8'h1C; mem['h1A63]=8'h46;
    mem['h1A64]=8'hAD; mem['h1A65]=8'h12; mem['h1A66]=8'h36; mem['h1A67]=8'h24;
    mem['h1A68]=8'h46; mem['h1A69]=8'hB6; mem['h1A6A]=8'h12; mem['h1A6B]=8'h46;
    mem['h1A6C]=8'h1A; mem['h1A6D]=8'h11; mem['h1A6E]=8'h36; mem['h1A6F]=8'h57;
    mem['h1A70]=8'hC7; mem['h1A71]=8'h3C; mem['h1A72]=8'hF7; mem['h1A73]=8'h44;
    mem['h1A74]=8'hF4; mem['h1A75]=8'h1A; mem['h1A76]=8'h36; mem['h1A77]=8'h1C;
    mem['h1A78]=8'hDD; mem['h1A79]=8'h26; mem['h1A7A]=8'h24; mem['h1A7B]=8'h0E;
    mem['h1A7C]=8'h04; mem['h1A7D]=8'h46; mem['h1A7E]=8'h0B; mem['h1A7F]=8'h11;
    mem['h1A80]=8'h44; mem['h1A81]=8'h47; mem['h1A82]=8'h1A; mem['h1A83]=8'h36;
    mem['h1A84]=8'h0B; mem['h1A85]=8'hC7; mem['h1A86]=8'h36; mem['h1A87]=8'h1F;
    mem['h1A88]=8'h87; mem['h1A89]=8'hF8; mem['h1A8A]=8'h36; mem['h1A8B]=8'h1C;
    mem['h1A8C]=8'h44; mem['h1A8D]=8'hA4; mem['h1A8E]=8'h12; mem['h1A8F]=8'h06;
    mem['h1A90]=8'hD3; mem['h1A91]=8'h16; mem['h1A92]=8'hD1; mem['h1A93]=8'h44;
    mem['h1A94]=8'h96; mem['h1A95]=8'h02; mem['h1A96]=8'hFF; mem['h1A97]=8'hFF;
    mem['h1A98]=8'hFF; mem['h1A99]=8'hFF; mem['h1A9A]=8'hFF; mem['h1A9B]=8'hFF;
    mem['h1A9C]=8'hFF; mem['h1A9D]=8'hFF; mem['h1A9E]=8'hFF; mem['h1A9F]=8'hFF;
    mem['h1AA0]=8'h36; mem['h1AA1]=8'h34; mem['h1AA2]=8'h2E; mem['h1AA3]=8'h01;
    mem['h1AA4]=8'h46; mem['h1AA5]=8'hA4; mem['h1AA6]=8'h12; mem['h1AA7]=8'h36;
    mem['h1AA8]=8'h28; mem['h1AA9]=8'h46; mem['h1AAA]=8'hB6; mem['h1AAB]=8'h12;
    mem['h1AAC]=8'h46; mem['h1AAD]=8'h26; mem['h1AAE]=8'h11; mem['h1AAF]=8'h36;
    mem['h1AB0]=8'h30; mem['h1AB1]=8'h46; mem['h1AB2]=8'hB6; mem['h1AB3]=8'h12;
    mem['h1AB4]=8'h46; mem['h1AB5]=8'h89; mem['h1AB6]=8'h10; mem['h1AB7]=8'h36;
    mem['h1AB8]=8'h34; mem['h1AB9]=8'h46; mem['h1ABA]=8'hAD; mem['h1ABB]=8'h12;
    mem['h1ABC]=8'h36; mem['h1ABD]=8'h57; mem['h1ABE]=8'hC7; mem['h1ABF]=8'h14;
    mem['h1AC0]=8'h10; mem['h1AC1]=8'hF8; mem['h1AC2]=8'h46; mem['h1AC3]=8'h00;
    mem['h1AC4]=8'h10; mem['h1AC5]=8'h36; mem['h1AC6]=8'h53; mem['h1AC7]=8'h3E;
    mem['h1AC8]=8'h00; mem['h1AC9]=8'h36; mem['h1ACA]=8'h57; mem['h1ACB]=8'h3E;
    mem['h1ACC]=8'h00; mem['h1ACD]=8'h46; mem['h1ACE]=8'h34; mem['h1ACF]=8'h10;
    mem['h1AD0]=8'h36; mem['h1AD1]=8'h57; mem['h1AD2]=8'hC7; mem['h1AD3]=8'h04;
    mem['h1AD4]=8'h10; mem['h1AD5]=8'hF8; mem['h1AD6]=8'h36; mem['h1AD7]=8'h34;
    mem['h1AD8]=8'h46; mem['h1AD9]=8'hB6; mem['h1ADA]=8'h12; mem['h1ADB]=8'h46;
    mem['h1ADC]=8'h1A; mem['h1ADD]=8'h11; mem['h1ADE]=8'h36; mem['h1ADF]=8'h34;
    mem['h1AE0]=8'h46; mem['h1AE1]=8'hAD; mem['h1AE2]=8'h12; mem['h1AE3]=8'h36;
    mem['h1AE4]=8'h57; mem['h1AE5]=8'hC7; mem['h1AE6]=8'h14; mem['h1AE7]=8'h10;
    mem['h1AE8]=8'hF8; mem['h1AE9]=8'h07; mem['h1AEA]=8'hFF; mem['h1AEB]=8'hFF;
    mem['h1AEC]=8'hFF; mem['h1AED]=8'hFF; mem['h1AEE]=8'hFF; mem['h1AEF]=8'hFF;
    mem['h1AF0]=8'hFF; mem['h1AF1]=8'hFF; mem['h1AF2]=8'hFF; mem['h1AF3]=8'hFF;
    mem['h1AF4]=8'h70; mem['h1AF5]=8'h83; mem['h1AF6]=8'h1A; mem['h1AF7]=8'h31;
    mem['h1AF8]=8'hC7; mem['h1AF9]=8'hA0; mem['h1AFA]=8'h68; mem['h1AFB]=8'h83;
    mem['h1AFC]=8'h1A; mem['h1AFD]=8'h44; mem['h1AFE]=8'h76; mem['h1AFF]=8'h1A;
    mem['h1B00]=8'hFF; mem['h1B01]=8'hFF; mem['h1B02]=8'hFF; mem['h1B03]=8'hFF;
    mem['h1B04]=8'hFF; mem['h1B05]=8'hFF; mem['h1B06]=8'hFF; mem['h1B07]=8'hFF;
    mem['h1B08]=8'hFF; mem['h1B09]=8'hFF; mem['h1B0A]=8'hFF; mem['h1B0B]=8'hFF;
    mem['h1B0C]=8'hFF; mem['h1B0D]=8'hFF; mem['h1B0E]=8'hFF; mem['h1B0F]=8'hFF;
    mem['h1B10]=8'hFF; mem['h1B11]=8'hFF; mem['h1B12]=8'hFF; mem['h1B13]=8'hFF;
    mem['h1B14]=8'hFF; mem['h1B15]=8'hFF; mem['h1B16]=8'hFF; mem['h1B17]=8'hFF;
    mem['h1B18]=8'hFF; mem['h1B19]=8'hFF; mem['h1B1A]=8'hFF; mem['h1B1B]=8'hFF;
    mem['h1B1C]=8'hFF; mem['h1B1D]=8'hFF; mem['h1B1E]=8'hFF; mem['h1B1F]=8'hFF;
    mem['h1B20]=8'hFF; mem['h1B21]=8'hFF; mem['h1B22]=8'hFF; mem['h1B23]=8'hFF;
    mem['h1B24]=8'hFF; mem['h1B25]=8'hFF; mem['h1B26]=8'hFF; mem['h1B27]=8'hFF;
    mem['h1B28]=8'hFF; mem['h1B29]=8'hFF; mem['h1B2A]=8'hFF; mem['h1B2B]=8'hFF;
    mem['h1B2C]=8'hFF; mem['h1B2D]=8'hFF; mem['h1B2E]=8'hFF; mem['h1B2F]=8'hFF;
    mem['h1B30]=8'hFF; mem['h1B31]=8'hFF; mem['h1B32]=8'hFF; mem['h1B33]=8'hFF;
    mem['h1B34]=8'hFF; mem['h1B35]=8'hFF; mem['h1B36]=8'hFF; mem['h1B37]=8'hFF;
    mem['h1B38]=8'hFF; mem['h1B39]=8'hFF; mem['h1B3A]=8'hFF; mem['h1B3B]=8'hFF;
    mem['h1B3C]=8'hFF; mem['h1B3D]=8'hFF; mem['h1B3E]=8'hFF; mem['h1B3F]=8'hFF;
    mem['h1B40]=8'hFF; mem['h1B41]=8'hFF; mem['h1B42]=8'hFF; mem['h1B43]=8'hFF;
    mem['h1B44]=8'hFF; mem['h1B45]=8'hFF; mem['h1B46]=8'hFF; mem['h1B47]=8'hFF;
    mem['h1B48]=8'hFF; mem['h1B49]=8'hFF; mem['h1B4A]=8'hFF; mem['h1B4B]=8'hFF;
    mem['h1B4C]=8'hFF; mem['h1B4D]=8'hFF; mem['h1B4E]=8'hFF; mem['h1B4F]=8'hFF;
    mem['h1B50]=8'hFF; mem['h1B51]=8'hFF; mem['h1B52]=8'hFF; mem['h1B53]=8'hFF;
    mem['h1B54]=8'hFF; mem['h1B55]=8'hFF; mem['h1B56]=8'hFF; mem['h1B57]=8'hFF;
    mem['h1B58]=8'hFF; mem['h1B59]=8'hFF; mem['h1B5A]=8'hFF; mem['h1B5B]=8'hFF;
    mem['h1B5C]=8'hFF; mem['h1B5D]=8'hFF; mem['h1B5E]=8'hFF; mem['h1B5F]=8'hFF;
    mem['h1B60]=8'hFF; mem['h1B61]=8'hFF; mem['h1B62]=8'hFF; mem['h1B63]=8'hFF;
    mem['h1B64]=8'hFF; mem['h1B65]=8'hFF; mem['h1B66]=8'hFF; mem['h1B67]=8'hFF;
    mem['h1B68]=8'hFF; mem['h1B69]=8'hFF; mem['h1B6A]=8'hFF; mem['h1B6B]=8'hFF;
    mem['h1B6C]=8'hFF; mem['h1B6D]=8'hFF; mem['h1B6E]=8'hFF; mem['h1B6F]=8'hFF;
    mem['h1B70]=8'hFF; mem['h1B71]=8'hFF; mem['h1B72]=8'hFF; mem['h1B73]=8'hFF;
    mem['h1B74]=8'hFF; mem['h1B75]=8'hFF; mem['h1B76]=8'hFF; mem['h1B77]=8'hFF;
    mem['h1B78]=8'hFF; mem['h1B79]=8'hFF; mem['h1B7A]=8'hFF; mem['h1B7B]=8'hFF;
    mem['h1B7C]=8'hFF; mem['h1B7D]=8'hFF; mem['h1B7E]=8'hFF; mem['h1B7F]=8'hFF;
    mem['h1B80]=8'hFF; mem['h1B81]=8'hFF; mem['h1B82]=8'hFF; mem['h1B83]=8'hFF;
    mem['h1B84]=8'hFF; mem['h1B85]=8'hFF; mem['h1B86]=8'hFF; mem['h1B87]=8'hFF;
    mem['h1B88]=8'hFF; mem['h1B89]=8'hFF; mem['h1B8A]=8'hFF; mem['h1B8B]=8'hFF;
    mem['h1B8C]=8'hFF; mem['h1B8D]=8'hFF; mem['h1B8E]=8'hFF; mem['h1B8F]=8'hFF;
    mem['h1B90]=8'hFF; mem['h1B91]=8'hFF; mem['h1B92]=8'hFF; mem['h1B93]=8'hFF;
    mem['h1B94]=8'hFF; mem['h1B95]=8'hFF; mem['h1B96]=8'hFF; mem['h1B97]=8'hFF;
    mem['h1B98]=8'hFF; mem['h1B99]=8'hFF; mem['h1B9A]=8'hFF; mem['h1B9B]=8'hFF;
    mem['h1B9C]=8'hFF; mem['h1B9D]=8'hFF; mem['h1B9E]=8'hFF; mem['h1B9F]=8'hFF;
    mem['h1BA0]=8'hFF; mem['h1BA1]=8'hFF; mem['h1BA2]=8'hFF; mem['h1BA3]=8'hFF;
    mem['h1BA4]=8'hFF; mem['h1BA5]=8'hFF; mem['h1BA6]=8'hFF; mem['h1BA7]=8'hFF;
    mem['h1BA8]=8'hFF; mem['h1BA9]=8'hFF; mem['h1BAA]=8'hFF; mem['h1BAB]=8'hFF;
    mem['h1BAC]=8'hFF; mem['h1BAD]=8'hFF; mem['h1BAE]=8'hFF; mem['h1BAF]=8'hFF;
    mem['h1BB0]=8'hFF; mem['h1BB1]=8'hFF; mem['h1BB2]=8'hFF; mem['h1BB3]=8'hFF;
    mem['h1BB4]=8'hFF; mem['h1BB5]=8'hFF; mem['h1BB6]=8'hFF; mem['h1BB7]=8'hFF;
    mem['h1BB8]=8'hFF; mem['h1BB9]=8'hFF; mem['h1BBA]=8'hFF; mem['h1BBB]=8'hFF;
    mem['h1BBC]=8'hFF; mem['h1BBD]=8'hFF; mem['h1BBE]=8'hFF; mem['h1BBF]=8'hFF;
    mem['h1BC0]=8'hFF; mem['h1BC1]=8'hFF; mem['h1BC2]=8'hFF; mem['h1BC3]=8'hFF;
    mem['h1BC4]=8'hFF; mem['h1BC5]=8'hFF; mem['h1BC6]=8'hFF; mem['h1BC7]=8'hFF;
    mem['h1BC8]=8'hFF; mem['h1BC9]=8'hFF; mem['h1BCA]=8'hFF; mem['h1BCB]=8'hFF;
    mem['h1BCC]=8'hFF; mem['h1BCD]=8'hFF; mem['h1BCE]=8'hFF; mem['h1BCF]=8'hFF;
    mem['h1BD0]=8'hFF; mem['h1BD1]=8'hFF; mem['h1BD2]=8'hFF; mem['h1BD3]=8'hFF;
    mem['h1BD4]=8'hFF; mem['h1BD5]=8'hFF; mem['h1BD6]=8'hFF; mem['h1BD7]=8'hFF;
    mem['h1BD8]=8'hFF; mem['h1BD9]=8'hFF; mem['h1BDA]=8'hFF; mem['h1BDB]=8'hFF;
    mem['h1BDC]=8'hFF; mem['h1BDD]=8'hFF; mem['h1BDE]=8'hFF; mem['h1BDF]=8'hFF;
    mem['h1BE0]=8'hFF; mem['h1BE1]=8'hFF; mem['h1BE2]=8'hFF; mem['h1BE3]=8'hFF;
    mem['h1BE4]=8'hFF; mem['h1BE5]=8'hFF; mem['h1BE6]=8'hFF; mem['h1BE7]=8'hFF;
    mem['h1BE8]=8'hFF; mem['h1BE9]=8'hFF; mem['h1BEA]=8'hFF; mem['h1BEB]=8'hFF;
    mem['h1BEC]=8'hFF; mem['h1BED]=8'hFF; mem['h1BEE]=8'hFF; mem['h1BEF]=8'hFF;
    mem['h1BF0]=8'hFF; mem['h1BF1]=8'hFF; mem['h1BF2]=8'hFF; mem['h1BF3]=8'hFF;
    mem['h1BF4]=8'hFF; mem['h1BF5]=8'hFF; mem['h1BF6]=8'hFF; mem['h1BF7]=8'hFF;
    mem['h1BF8]=8'hFF; mem['h1BF9]=8'hFF; mem['h1BFA]=8'hFF; mem['h1BFB]=8'hFF;
    mem['h1BFC]=8'hFF; mem['h1BFD]=8'hFF; mem['h1BFE]=8'hFF; mem['h1BFF]=8'hFF;
    mem['h1C00]=8'hFF; mem['h1C01]=8'hFF; mem['h1C02]=8'hFF; mem['h1C03]=8'hFF;
    mem['h1C04]=8'hFF; mem['h1C05]=8'hFF; mem['h1C06]=8'hFF; mem['h1C07]=8'hFF;
    mem['h1C08]=8'hFF; mem['h1C09]=8'hFF; mem['h1C0A]=8'hFF; mem['h1C0B]=8'hFF;
    mem['h1C0C]=8'hFF; mem['h1C0D]=8'hFF; mem['h1C0E]=8'hFF; mem['h1C0F]=8'hFF;
    mem['h1C10]=8'hFF; mem['h1C11]=8'hFF; mem['h1C12]=8'hFF; mem['h1C13]=8'hFF;
    mem['h1C14]=8'hFF; mem['h1C15]=8'hFF; mem['h1C16]=8'hFF; mem['h1C17]=8'hFF;
    mem['h1C18]=8'hFF; mem['h1C19]=8'hFF; mem['h1C1A]=8'hFF; mem['h1C1B]=8'hFF;
    mem['h1C1C]=8'hFF; mem['h1C1D]=8'hFF; mem['h1C1E]=8'hFF; mem['h1C1F]=8'hFF;
    mem['h1C20]=8'hFF; mem['h1C21]=8'hFF; mem['h1C22]=8'hFF; mem['h1C23]=8'hFF;
    mem['h1C24]=8'hFF; mem['h1C25]=8'hFF; mem['h1C26]=8'hFF; mem['h1C27]=8'hFF;
    mem['h1C28]=8'hFF; mem['h1C29]=8'hFF; mem['h1C2A]=8'hFF; mem['h1C2B]=8'hFF;
    mem['h1C2C]=8'hFF; mem['h1C2D]=8'hFF; mem['h1C2E]=8'hFF; mem['h1C2F]=8'hFF;
    mem['h1C30]=8'hFF; mem['h1C31]=8'hFF; mem['h1C32]=8'hFF; mem['h1C33]=8'hFF;
    mem['h1C34]=8'hFF; mem['h1C35]=8'hFF; mem['h1C36]=8'hFF; mem['h1C37]=8'hFF;
    mem['h1C38]=8'hFF; mem['h1C39]=8'hFF; mem['h1C3A]=8'hFF; mem['h1C3B]=8'hFF;
    mem['h1C3C]=8'hFF; mem['h1C3D]=8'hFF; mem['h1C3E]=8'hFF; mem['h1C3F]=8'hFF;
    mem['h1C40]=8'hFF; mem['h1C41]=8'hFF; mem['h1C42]=8'hFF; mem['h1C43]=8'hFF;
    mem['h1C44]=8'hFF; mem['h1C45]=8'hFF; mem['h1C46]=8'hFF; mem['h1C47]=8'hFF;
    mem['h1C48]=8'hFF; mem['h1C49]=8'hFF; mem['h1C4A]=8'hFF; mem['h1C4B]=8'hFF;
    mem['h1C4C]=8'hFF; mem['h1C4D]=8'hFF; mem['h1C4E]=8'hFF; mem['h1C4F]=8'hFF;
    mem['h1C50]=8'hFF; mem['h1C51]=8'hFF; mem['h1C52]=8'hFF; mem['h1C53]=8'hFF;
    mem['h1C54]=8'hFF; mem['h1C55]=8'hFF; mem['h1C56]=8'hFF; mem['h1C57]=8'hFF;
    mem['h1C58]=8'hFF; mem['h1C59]=8'hFF; mem['h1C5A]=8'hFF; mem['h1C5B]=8'hFF;
    mem['h1C5C]=8'hFF; mem['h1C5D]=8'hFF; mem['h1C5E]=8'hFF; mem['h1C5F]=8'hFF;
    mem['h1C60]=8'hFF; mem['h1C61]=8'hFF; mem['h1C62]=8'hFF; mem['h1C63]=8'hFF;
    mem['h1C64]=8'hFF; mem['h1C65]=8'hFF; mem['h1C66]=8'hFF; mem['h1C67]=8'hFF;
    mem['h1C68]=8'hFF; mem['h1C69]=8'hFF; mem['h1C6A]=8'hFF; mem['h1C6B]=8'hFF;
    mem['h1C6C]=8'hFF; mem['h1C6D]=8'hFF; mem['h1C6E]=8'hFF; mem['h1C6F]=8'hFF;
    mem['h1C70]=8'hFF; mem['h1C71]=8'hFF; mem['h1C72]=8'hFF; mem['h1C73]=8'hFF;
    mem['h1C74]=8'hFF; mem['h1C75]=8'hFF; mem['h1C76]=8'hFF; mem['h1C77]=8'hFF;
    mem['h1C78]=8'hFF; mem['h1C79]=8'hFF; mem['h1C7A]=8'hFF; mem['h1C7B]=8'hFF;
    mem['h1C7C]=8'hFF; mem['h1C7D]=8'hFF; mem['h1C7E]=8'hFF; mem['h1C7F]=8'hFF;
    mem['h1C80]=8'hFF; mem['h1C81]=8'hFF; mem['h1C82]=8'hFF; mem['h1C83]=8'hFF;
    mem['h1C84]=8'hFF; mem['h1C85]=8'hFF; mem['h1C86]=8'hFF; mem['h1C87]=8'hFF;
    mem['h1C88]=8'hFF; mem['h1C89]=8'hFF; mem['h1C8A]=8'hFF; mem['h1C8B]=8'hFF;
    mem['h1C8C]=8'hFF; mem['h1C8D]=8'hFF; mem['h1C8E]=8'hFF; mem['h1C8F]=8'hFF;
    mem['h1C90]=8'hFF; mem['h1C91]=8'hFF; mem['h1C92]=8'hFF; mem['h1C93]=8'hFF;
    mem['h1C94]=8'hFF; mem['h1C95]=8'hFF; mem['h1C96]=8'hFF; mem['h1C97]=8'hFF;
    mem['h1C98]=8'hFF; mem['h1C99]=8'hFF; mem['h1C9A]=8'hFF; mem['h1C9B]=8'hFF;
    mem['h1C9C]=8'hFF; mem['h1C9D]=8'hFF; mem['h1C9E]=8'hFF; mem['h1C9F]=8'hFF;
    mem['h1CA0]=8'hFF; mem['h1CA1]=8'hFF; mem['h1CA2]=8'hFF; mem['h1CA3]=8'hFF;
    mem['h1CA4]=8'hFF; mem['h1CA5]=8'hFF; mem['h1CA6]=8'hFF; mem['h1CA7]=8'hFF;
    mem['h1CA8]=8'hFF; mem['h1CA9]=8'hFF; mem['h1CAA]=8'hFF; mem['h1CAB]=8'hFF;
    mem['h1CAC]=8'hFF; mem['h1CAD]=8'hFF; mem['h1CAE]=8'hFF; mem['h1CAF]=8'hFF;
    mem['h1CB0]=8'hFF; mem['h1CB1]=8'hFF; mem['h1CB2]=8'hFF; mem['h1CB3]=8'hFF;
    mem['h1CB4]=8'hFF; mem['h1CB5]=8'hFF; mem['h1CB6]=8'hFF; mem['h1CB7]=8'hFF;
    mem['h1CB8]=8'hFF; mem['h1CB9]=8'hFF; mem['h1CBA]=8'hFF; mem['h1CBB]=8'hFF;
    mem['h1CBC]=8'hFF; mem['h1CBD]=8'hFF; mem['h1CBE]=8'hFF; mem['h1CBF]=8'hFF;
    mem['h1CC0]=8'hFF; mem['h1CC1]=8'hFF; mem['h1CC2]=8'hFF; mem['h1CC3]=8'hFF;
    mem['h1CC4]=8'hFF; mem['h1CC5]=8'hFF; mem['h1CC6]=8'hFF; mem['h1CC7]=8'hFF;
    mem['h1CC8]=8'hFF; mem['h1CC9]=8'hFF; mem['h1CCA]=8'hFF; mem['h1CCB]=8'hFF;
    mem['h1CCC]=8'hFF; mem['h1CCD]=8'hFF; mem['h1CCE]=8'hFF; mem['h1CCF]=8'hFF;
    mem['h1CD0]=8'hFF; mem['h1CD1]=8'hFF; mem['h1CD2]=8'hFF; mem['h1CD3]=8'hFF;
    mem['h1CD4]=8'hFF; mem['h1CD5]=8'hFF; mem['h1CD6]=8'hFF; mem['h1CD7]=8'hFF;
    mem['h1CD8]=8'hFF; mem['h1CD9]=8'hFF; mem['h1CDA]=8'hFF; mem['h1CDB]=8'hFF;
    mem['h1CDC]=8'hFF; mem['h1CDD]=8'hFF; mem['h1CDE]=8'hFF; mem['h1CDF]=8'hFF;
    mem['h1CE0]=8'hFF; mem['h1CE1]=8'hFF; mem['h1CE2]=8'hFF; mem['h1CE3]=8'hFF;
    mem['h1CE4]=8'hFF; mem['h1CE5]=8'hFF; mem['h1CE6]=8'hFF; mem['h1CE7]=8'hFF;
    mem['h1CE8]=8'hFF; mem['h1CE9]=8'hFF; mem['h1CEA]=8'hFF; mem['h1CEB]=8'hFF;
    mem['h1CEC]=8'hFF; mem['h1CED]=8'hFF; mem['h1CEE]=8'hFF; mem['h1CEF]=8'hFF;
    mem['h1CF0]=8'hFF; mem['h1CF1]=8'hFF; mem['h1CF2]=8'hFF; mem['h1CF3]=8'hFF;
    mem['h1CF4]=8'hFF; mem['h1CF5]=8'hFF; mem['h1CF6]=8'hFF; mem['h1CF7]=8'hFF;
    mem['h1CF8]=8'hFF; mem['h1CF9]=8'hFF; mem['h1CFA]=8'hFF; mem['h1CFB]=8'hFF;
    mem['h1CFC]=8'hFF; mem['h1CFD]=8'hFF; mem['h1CFE]=8'hFF; mem['h1CFF]=8'hFF;
    mem['h1D00]=8'hFF; mem['h1D01]=8'hFF; mem['h1D02]=8'hFF; mem['h1D03]=8'hFF;
    mem['h1D04]=8'hFF; mem['h1D05]=8'hFF; mem['h1D06]=8'hFF; mem['h1D07]=8'hFF;
    mem['h1D08]=8'hFF; mem['h1D09]=8'hFF; mem['h1D0A]=8'hFF; mem['h1D0B]=8'hFF;
    mem['h1D0C]=8'hFF; mem['h1D0D]=8'hFF; mem['h1D0E]=8'hFF; mem['h1D0F]=8'hFF;
    mem['h1D10]=8'hFF; mem['h1D11]=8'hFF; mem['h1D12]=8'hFF; mem['h1D13]=8'hFF;
    mem['h1D14]=8'hFF; mem['h1D15]=8'hFF; mem['h1D16]=8'hFF; mem['h1D17]=8'hFF;
    mem['h1D18]=8'hFF; mem['h1D19]=8'hFF; mem['h1D1A]=8'hFF; mem['h1D1B]=8'hFF;
    mem['h1D1C]=8'hFF; mem['h1D1D]=8'hFF; mem['h1D1E]=8'hFF; mem['h1D1F]=8'hFF;
    mem['h1D20]=8'hFF; mem['h1D21]=8'hFF; mem['h1D22]=8'hFF; mem['h1D23]=8'hFF;
    mem['h1D24]=8'hFF; mem['h1D25]=8'hFF; mem['h1D26]=8'hFF; mem['h1D27]=8'hFF;
    mem['h1D28]=8'hFF; mem['h1D29]=8'hFF; mem['h1D2A]=8'hFF; mem['h1D2B]=8'hFF;
    mem['h1D2C]=8'hFF; mem['h1D2D]=8'hFF; mem['h1D2E]=8'hFF; mem['h1D2F]=8'hFF;
    mem['h1D30]=8'hFF; mem['h1D31]=8'hFF; mem['h1D32]=8'hFF; mem['h1D33]=8'hFF;
    mem['h1D34]=8'hFF; mem['h1D35]=8'hFF; mem['h1D36]=8'hFF; mem['h1D37]=8'hFF;
    mem['h1D38]=8'hFF; mem['h1D39]=8'hFF; mem['h1D3A]=8'hFF; mem['h1D3B]=8'hFF;
    mem['h1D3C]=8'hFF; mem['h1D3D]=8'hFF; mem['h1D3E]=8'hFF; mem['h1D3F]=8'hFF;
    mem['h1D40]=8'hFF; mem['h1D41]=8'hFF; mem['h1D42]=8'hFF; mem['h1D43]=8'hFF;
    mem['h1D44]=8'hFF; mem['h1D45]=8'hFF; mem['h1D46]=8'hFF; mem['h1D47]=8'hFF;
    mem['h1D48]=8'hFF; mem['h1D49]=8'hFF; mem['h1D4A]=8'hFF; mem['h1D4B]=8'hFF;
    mem['h1D4C]=8'hFF; mem['h1D4D]=8'hFF; mem['h1D4E]=8'hFF; mem['h1D4F]=8'hFF;
    mem['h1D50]=8'hFF; mem['h1D51]=8'hFF; mem['h1D52]=8'hFF; mem['h1D53]=8'hFF;
    mem['h1D54]=8'hFF; mem['h1D55]=8'hFF; mem['h1D56]=8'hFF; mem['h1D57]=8'hFF;
    mem['h1D58]=8'hFF; mem['h1D59]=8'hFF; mem['h1D5A]=8'hFF; mem['h1D5B]=8'hFF;
    mem['h1D5C]=8'hFF; mem['h1D5D]=8'hFF; mem['h1D5E]=8'hFF; mem['h1D5F]=8'hFF;
    mem['h1D60]=8'hFF; mem['h1D61]=8'hFF; mem['h1D62]=8'hFF; mem['h1D63]=8'hFF;
    mem['h1D64]=8'hFF; mem['h1D65]=8'hFF; mem['h1D66]=8'hFF; mem['h1D67]=8'hFF;
    mem['h1D68]=8'hFF; mem['h1D69]=8'hFF; mem['h1D6A]=8'hFF; mem['h1D6B]=8'hFF;
    mem['h1D6C]=8'hFF; mem['h1D6D]=8'hFF; mem['h1D6E]=8'hFF; mem['h1D6F]=8'hFF;
    mem['h1D70]=8'hFF; mem['h1D71]=8'hFF; mem['h1D72]=8'hFF; mem['h1D73]=8'hFF;
    mem['h1D74]=8'hFF; mem['h1D75]=8'hFF; mem['h1D76]=8'hFF; mem['h1D77]=8'hFF;
    mem['h1D78]=8'hFF; mem['h1D79]=8'hFF; mem['h1D7A]=8'hFF; mem['h1D7B]=8'hFF;
    mem['h1D7C]=8'hFF; mem['h1D7D]=8'hFF; mem['h1D7E]=8'hFF; mem['h1D7F]=8'hFF;
    mem['h1D80]=8'hFF; mem['h1D81]=8'hFF; mem['h1D82]=8'hFF; mem['h1D83]=8'hFF;
    mem['h1D84]=8'hFF; mem['h1D85]=8'hFF; mem['h1D86]=8'hFF; mem['h1D87]=8'hFF;
    mem['h1D88]=8'hFF; mem['h1D89]=8'hFF; mem['h1D8A]=8'hFF; mem['h1D8B]=8'hFF;
    mem['h1D8C]=8'hFF; mem['h1D8D]=8'hFF; mem['h1D8E]=8'hFF; mem['h1D8F]=8'hFF;
    mem['h1D90]=8'hFF; mem['h1D91]=8'hFF; mem['h1D92]=8'hFF; mem['h1D93]=8'hFF;
    mem['h1D94]=8'hFF; mem['h1D95]=8'hFF; mem['h1D96]=8'hFF; mem['h1D97]=8'hFF;
    mem['h1D98]=8'hFF; mem['h1D99]=8'hFF; mem['h1D9A]=8'hFF; mem['h1D9B]=8'hFF;
    mem['h1D9C]=8'hFF; mem['h1D9D]=8'hFF; mem['h1D9E]=8'hFF; mem['h1D9F]=8'hFF;
    mem['h1DA0]=8'hFF; mem['h1DA1]=8'hFF; mem['h1DA2]=8'hFF; mem['h1DA3]=8'hFF;
    mem['h1DA4]=8'hFF; mem['h1DA5]=8'hFF; mem['h1DA6]=8'hFF; mem['h1DA7]=8'hFF;
    mem['h1DA8]=8'hFF; mem['h1DA9]=8'hFF; mem['h1DAA]=8'hFF; mem['h1DAB]=8'hFF;
    mem['h1DAC]=8'hFF; mem['h1DAD]=8'hFF; mem['h1DAE]=8'hFF; mem['h1DAF]=8'hFF;
    mem['h1DB0]=8'hFF; mem['h1DB1]=8'hFF; mem['h1DB2]=8'hFF; mem['h1DB3]=8'hFF;
    mem['h1DB4]=8'hFF; mem['h1DB5]=8'hFF; mem['h1DB6]=8'hFF; mem['h1DB7]=8'hFF;
    mem['h1DB8]=8'hFF; mem['h1DB9]=8'hFF; mem['h1DBA]=8'hFF; mem['h1DBB]=8'hFF;
    mem['h1DBC]=8'hFF; mem['h1DBD]=8'hFF; mem['h1DBE]=8'hFF; mem['h1DBF]=8'hFF;
    mem['h1DC0]=8'hFF; mem['h1DC1]=8'hFF; mem['h1DC2]=8'hFF; mem['h1DC3]=8'hFF;
    mem['h1DC4]=8'hFF; mem['h1DC5]=8'hFF; mem['h1DC6]=8'hFF; mem['h1DC7]=8'hFF;
    mem['h1DC8]=8'hFF; mem['h1DC9]=8'hFF; mem['h1DCA]=8'hFF; mem['h1DCB]=8'hFF;
    mem['h1DCC]=8'hFF; mem['h1DCD]=8'hFF; mem['h1DCE]=8'hFF; mem['h1DCF]=8'hFF;
    mem['h1DD0]=8'hFF; mem['h1DD1]=8'hFF; mem['h1DD2]=8'hFF; mem['h1DD3]=8'hFF;
    mem['h1DD4]=8'hFF; mem['h1DD5]=8'hFF; mem['h1DD6]=8'hFF; mem['h1DD7]=8'hFF;
    mem['h1DD8]=8'hFF; mem['h1DD9]=8'hFF; mem['h1DDA]=8'hFF; mem['h1DDB]=8'hFF;
    mem['h1DDC]=8'hFF; mem['h1DDD]=8'hFF; mem['h1DDE]=8'hFF; mem['h1DDF]=8'hFF;
    mem['h1DE0]=8'hFF; mem['h1DE1]=8'hFF; mem['h1DE2]=8'hFF; mem['h1DE3]=8'hFF;
    mem['h1DE4]=8'hFF; mem['h1DE5]=8'hFF; mem['h1DE6]=8'hFF; mem['h1DE7]=8'hFF;
    mem['h1DE8]=8'hFF; mem['h1DE9]=8'hFF; mem['h1DEA]=8'hFF; mem['h1DEB]=8'hFF;
    mem['h1DEC]=8'hFF; mem['h1DED]=8'hFF; mem['h1DEE]=8'hFF; mem['h1DEF]=8'hFF;
    mem['h1DF0]=8'hFF; mem['h1DF1]=8'hFF; mem['h1DF2]=8'hFF; mem['h1DF3]=8'hFF;
    mem['h1DF4]=8'hFF; mem['h1DF5]=8'hFF; mem['h1DF6]=8'hFF; mem['h1DF7]=8'hFF;
    mem['h1DF8]=8'hFF; mem['h1DF9]=8'hFF; mem['h1DFA]=8'hFF; mem['h1DFB]=8'hFF;
    mem['h1DFC]=8'hFF; mem['h1DFD]=8'hFF; mem['h1DFE]=8'hFF; mem['h1DFF]=8'hFF;
    mem['h1E00]=8'hFF; mem['h1E01]=8'hFF; mem['h1E02]=8'hFF; mem['h1E03]=8'hFF;
    mem['h1E04]=8'hFF; mem['h1E05]=8'hFF; mem['h1E06]=8'hFF; mem['h1E07]=8'hFF;
    mem['h1E08]=8'hFF; mem['h1E09]=8'hFF; mem['h1E0A]=8'hFF; mem['h1E0B]=8'hFF;
    mem['h1E0C]=8'hFF; mem['h1E0D]=8'hFF; mem['h1E0E]=8'hFF; mem['h1E0F]=8'hFF;
    mem['h1E10]=8'hFF; mem['h1E11]=8'hFF; mem['h1E12]=8'hFF; mem['h1E13]=8'hFF;
    mem['h1E14]=8'hFF; mem['h1E15]=8'hFF; mem['h1E16]=8'hFF; mem['h1E17]=8'hFF;
    mem['h1E18]=8'hFF; mem['h1E19]=8'hFF; mem['h1E1A]=8'hFF; mem['h1E1B]=8'hFF;
    mem['h1E1C]=8'hFF; mem['h1E1D]=8'hFF; mem['h1E1E]=8'hFF; mem['h1E1F]=8'hFF;
    mem['h1E20]=8'hFF; mem['h1E21]=8'hFF; mem['h1E22]=8'hFF; mem['h1E23]=8'hFF;
    mem['h1E24]=8'hFF; mem['h1E25]=8'hFF; mem['h1E26]=8'hFF; mem['h1E27]=8'hFF;
    mem['h1E28]=8'hFF; mem['h1E29]=8'hFF; mem['h1E2A]=8'hFF; mem['h1E2B]=8'hFF;
    mem['h1E2C]=8'hFF; mem['h1E2D]=8'hFF; mem['h1E2E]=8'hFF; mem['h1E2F]=8'hFF;
    mem['h1E30]=8'hFF; mem['h1E31]=8'hFF; mem['h1E32]=8'hFF; mem['h1E33]=8'hFF;
    mem['h1E34]=8'hFF; mem['h1E35]=8'hFF; mem['h1E36]=8'hFF; mem['h1E37]=8'hFF;
    mem['h1E38]=8'hFF; mem['h1E39]=8'hFF; mem['h1E3A]=8'hFF; mem['h1E3B]=8'hFF;
    mem['h1E3C]=8'hFF; mem['h1E3D]=8'hFF; mem['h1E3E]=8'hFF; mem['h1E3F]=8'hFF;
    mem['h1E40]=8'hFF; mem['h1E41]=8'hFF; mem['h1E42]=8'hFF; mem['h1E43]=8'hFF;
    mem['h1E44]=8'hFF; mem['h1E45]=8'hFF; mem['h1E46]=8'hFF; mem['h1E47]=8'hFF;
    mem['h1E48]=8'hFF; mem['h1E49]=8'hFF; mem['h1E4A]=8'hFF; mem['h1E4B]=8'hFF;
    mem['h1E4C]=8'hFF; mem['h1E4D]=8'hFF; mem['h1E4E]=8'hFF; mem['h1E4F]=8'hFF;
    mem['h1E50]=8'hFF; mem['h1E51]=8'hFF; mem['h1E52]=8'hFF; mem['h1E53]=8'hFF;
    mem['h1E54]=8'hFF; mem['h1E55]=8'hFF; mem['h1E56]=8'hFF; mem['h1E57]=8'hFF;
    mem['h1E58]=8'hFF; mem['h1E59]=8'hFF; mem['h1E5A]=8'hFF; mem['h1E5B]=8'hFF;
    mem['h1E5C]=8'hFF; mem['h1E5D]=8'hFF; mem['h1E5E]=8'hFF; mem['h1E5F]=8'hFF;
    mem['h1E60]=8'hFF; mem['h1E61]=8'hFF; mem['h1E62]=8'hFF; mem['h1E63]=8'hFF;
    mem['h1E64]=8'hFF; mem['h1E65]=8'hFF; mem['h1E66]=8'hFF; mem['h1E67]=8'hFF;
    mem['h1E68]=8'hFF; mem['h1E69]=8'hFF; mem['h1E6A]=8'hFF; mem['h1E6B]=8'hFF;
    mem['h1E6C]=8'hFF; mem['h1E6D]=8'hFF; mem['h1E6E]=8'hFF; mem['h1E6F]=8'hFF;
    mem['h1E70]=8'hFF; mem['h1E71]=8'hFF; mem['h1E72]=8'hFF; mem['h1E73]=8'hFF;
    mem['h1E74]=8'hFF; mem['h1E75]=8'hFF; mem['h1E76]=8'hFF; mem['h1E77]=8'hFF;
    mem['h1E78]=8'hFF; mem['h1E79]=8'hFF; mem['h1E7A]=8'hFF; mem['h1E7B]=8'hFF;
    mem['h1E7C]=8'hFF; mem['h1E7D]=8'hFF; mem['h1E7E]=8'hFF; mem['h1E7F]=8'hFF;
    mem['h1E80]=8'hFF; mem['h1E81]=8'hFF; mem['h1E82]=8'hFF; mem['h1E83]=8'hFF;
    mem['h1E84]=8'hFF; mem['h1E85]=8'hFF; mem['h1E86]=8'hFF; mem['h1E87]=8'hFF;
    mem['h1E88]=8'hFF; mem['h1E89]=8'hFF; mem['h1E8A]=8'hFF; mem['h1E8B]=8'hFF;
    mem['h1E8C]=8'hFF; mem['h1E8D]=8'hFF; mem['h1E8E]=8'hFF; mem['h1E8F]=8'hFF;
    mem['h1E90]=8'hFF; mem['h1E91]=8'hFF; mem['h1E92]=8'hFF; mem['h1E93]=8'hFF;
    mem['h1E94]=8'hFF; mem['h1E95]=8'hFF; mem['h1E96]=8'hFF; mem['h1E97]=8'hFF;
    mem['h1E98]=8'hFF; mem['h1E99]=8'hFF; mem['h1E9A]=8'hFF; mem['h1E9B]=8'hFF;
    mem['h1E9C]=8'hFF; mem['h1E9D]=8'hFF; mem['h1E9E]=8'hFF; mem['h1E9F]=8'hFF;
    mem['h1EA0]=8'hFF; mem['h1EA1]=8'hFF; mem['h1EA2]=8'hFF; mem['h1EA3]=8'hFF;
    mem['h1EA4]=8'hFF; mem['h1EA5]=8'hFF; mem['h1EA6]=8'hFF; mem['h1EA7]=8'hFF;
    mem['h1EA8]=8'hFF; mem['h1EA9]=8'hFF; mem['h1EAA]=8'hFF; mem['h1EAB]=8'hFF;
    mem['h1EAC]=8'hFF; mem['h1EAD]=8'hFF; mem['h1EAE]=8'hFF; mem['h1EAF]=8'hFF;
    mem['h1EB0]=8'hFF; mem['h1EB1]=8'hFF; mem['h1EB2]=8'hFF; mem['h1EB3]=8'hFF;
    mem['h1EB4]=8'hFF; mem['h1EB5]=8'hFF; mem['h1EB6]=8'hFF; mem['h1EB7]=8'hFF;
    mem['h1EB8]=8'hFF; mem['h1EB9]=8'hFF; mem['h1EBA]=8'hFF; mem['h1EBB]=8'hFF;
    mem['h1EBC]=8'hFF; mem['h1EBD]=8'hFF; mem['h1EBE]=8'hFF; mem['h1EBF]=8'hFF;
    mem['h1EC0]=8'hFF; mem['h1EC1]=8'hFF; mem['h1EC2]=8'hFF; mem['h1EC3]=8'hFF;
    mem['h1EC4]=8'hFF; mem['h1EC5]=8'hFF; mem['h1EC6]=8'hFF; mem['h1EC7]=8'hFF;
    mem['h1EC8]=8'hFF; mem['h1EC9]=8'hFF; mem['h1ECA]=8'hFF; mem['h1ECB]=8'hFF;
    mem['h1ECC]=8'hFF; mem['h1ECD]=8'hFF; mem['h1ECE]=8'hFF; mem['h1ECF]=8'hFF;
    mem['h1ED0]=8'hFF; mem['h1ED1]=8'hFF; mem['h1ED2]=8'hFF; mem['h1ED3]=8'hFF;
    mem['h1ED4]=8'hFF; mem['h1ED5]=8'hFF; mem['h1ED6]=8'hFF; mem['h1ED7]=8'hFF;
    mem['h1ED8]=8'hFF; mem['h1ED9]=8'hFF; mem['h1EDA]=8'hFF; mem['h1EDB]=8'hFF;
    mem['h1EDC]=8'hFF; mem['h1EDD]=8'hFF; mem['h1EDE]=8'hFF; mem['h1EDF]=8'hFF;
    mem['h1EE0]=8'hFF; mem['h1EE1]=8'hFF; mem['h1EE2]=8'hFF; mem['h1EE3]=8'hFF;
    mem['h1EE4]=8'hFF; mem['h1EE5]=8'hFF; mem['h1EE6]=8'hFF; mem['h1EE7]=8'hFF;
    mem['h1EE8]=8'hFF; mem['h1EE9]=8'hFF; mem['h1EEA]=8'hFF; mem['h1EEB]=8'hFF;
    mem['h1EEC]=8'hFF; mem['h1EED]=8'hFF; mem['h1EEE]=8'hFF; mem['h1EEF]=8'hFF;
    mem['h1EF0]=8'hFF; mem['h1EF1]=8'hFF; mem['h1EF2]=8'hFF; mem['h1EF3]=8'hFF;
    mem['h1EF4]=8'hFF; mem['h1EF5]=8'hFF; mem['h1EF6]=8'hFF; mem['h1EF7]=8'hFF;
    mem['h1EF8]=8'hFF; mem['h1EF9]=8'hFF; mem['h1EFA]=8'hFF; mem['h1EFB]=8'hFF;
    mem['h1EFC]=8'hFF; mem['h1EFD]=8'hFF; mem['h1EFE]=8'hFF; mem['h1EFF]=8'hFF;
    mem['h1F00]=8'hFF; mem['h1F01]=8'hFF; mem['h1F02]=8'hFF; mem['h1F03]=8'hFF;
    mem['h1F04]=8'hFF; mem['h1F05]=8'hFF; mem['h1F06]=8'hFF; mem['h1F07]=8'hFF;
    mem['h1F08]=8'hFF; mem['h1F09]=8'hFF; mem['h1F0A]=8'hFF; mem['h1F0B]=8'hFF;
    mem['h1F0C]=8'hFF; mem['h1F0D]=8'hFF; mem['h1F0E]=8'hFF; mem['h1F0F]=8'hFF;
    mem['h1F10]=8'hFF; mem['h1F11]=8'hFF; mem['h1F12]=8'hFF; mem['h1F13]=8'hFF;
    mem['h1F14]=8'hFF; mem['h1F15]=8'hFF; mem['h1F16]=8'hFF; mem['h1F17]=8'hFF;
    mem['h1F18]=8'hFF; mem['h1F19]=8'hFF; mem['h1F1A]=8'hFF; mem['h1F1B]=8'hFF;
    mem['h1F1C]=8'hFF; mem['h1F1D]=8'hFF; mem['h1F1E]=8'hFF; mem['h1F1F]=8'hFF;
    mem['h1F20]=8'hFF; mem['h1F21]=8'hFF; mem['h1F22]=8'hFF; mem['h1F23]=8'hFF;
    mem['h1F24]=8'hFF; mem['h1F25]=8'hFF; mem['h1F26]=8'hFF; mem['h1F27]=8'hFF;
    mem['h1F28]=8'hFF; mem['h1F29]=8'hFF; mem['h1F2A]=8'hFF; mem['h1F2B]=8'hFF;
    mem['h1F2C]=8'hFF; mem['h1F2D]=8'hFF; mem['h1F2E]=8'hFF; mem['h1F2F]=8'hFF;
    mem['h1F30]=8'hFF; mem['h1F31]=8'hFF; mem['h1F32]=8'hFF; mem['h1F33]=8'hFF;
    mem['h1F34]=8'hFF; mem['h1F35]=8'hFF; mem['h1F36]=8'hFF; mem['h1F37]=8'hFF;
    mem['h1F38]=8'hFF; mem['h1F39]=8'hFF; mem['h1F3A]=8'hFF; mem['h1F3B]=8'hFF;
    mem['h1F3C]=8'hFF; mem['h1F3D]=8'hFF; mem['h1F3E]=8'hFF; mem['h1F3F]=8'hFF;
    mem['h1F40]=8'hFF; mem['h1F41]=8'hFF; mem['h1F42]=8'hFF; mem['h1F43]=8'hFF;
    mem['h1F44]=8'hFF; mem['h1F45]=8'hFF; mem['h1F46]=8'hFF; mem['h1F47]=8'hFF;
    mem['h1F48]=8'hFF; mem['h1F49]=8'hFF; mem['h1F4A]=8'hFF; mem['h1F4B]=8'hFF;
    mem['h1F4C]=8'hFF; mem['h1F4D]=8'hFF; mem['h1F4E]=8'hFF; mem['h1F4F]=8'hFF;
    mem['h1F50]=8'hFF; mem['h1F51]=8'hFF; mem['h1F52]=8'hFF; mem['h1F53]=8'hFF;
    mem['h1F54]=8'hFF; mem['h1F55]=8'hFF; mem['h1F56]=8'hFF; mem['h1F57]=8'hFF;
    mem['h1F58]=8'hFF; mem['h1F59]=8'hFF; mem['h1F5A]=8'hFF; mem['h1F5B]=8'hFF;
    mem['h1F5C]=8'hFF; mem['h1F5D]=8'hFF; mem['h1F5E]=8'hFF; mem['h1F5F]=8'hFF;
    mem['h1F60]=8'hFF; mem['h1F61]=8'hFF; mem['h1F62]=8'hFF; mem['h1F63]=8'hFF;
    mem['h1F64]=8'hFF; mem['h1F65]=8'hFF; mem['h1F66]=8'hFF; mem['h1F67]=8'hFF;
    mem['h1F68]=8'hFF; mem['h1F69]=8'hFF; mem['h1F6A]=8'hFF; mem['h1F6B]=8'hFF;
    mem['h1F6C]=8'hFF; mem['h1F6D]=8'hFF; mem['h1F6E]=8'hFF; mem['h1F6F]=8'hFF;
    mem['h1F70]=8'hFF; mem['h1F71]=8'hFF; mem['h1F72]=8'hFF; mem['h1F73]=8'hFF;
    mem['h1F74]=8'hFF; mem['h1F75]=8'hFF; mem['h1F76]=8'hFF; mem['h1F77]=8'hFF;
    mem['h1F78]=8'hFF; mem['h1F79]=8'hFF; mem['h1F7A]=8'hFF; mem['h1F7B]=8'hFF;
    mem['h1F7C]=8'hFF; mem['h1F7D]=8'hFF; mem['h1F7E]=8'hFF; mem['h1F7F]=8'hFF;
    mem['h1F80]=8'hFF; mem['h1F81]=8'hFF; mem['h1F82]=8'hFF; mem['h1F83]=8'hFF;
    mem['h1F84]=8'hFF; mem['h1F85]=8'hFF; mem['h1F86]=8'hFF; mem['h1F87]=8'hFF;
    mem['h1F88]=8'hFF; mem['h1F89]=8'hFF; mem['h1F8A]=8'hFF; mem['h1F8B]=8'hFF;
    mem['h1F8C]=8'hFF; mem['h1F8D]=8'hFF; mem['h1F8E]=8'hFF; mem['h1F8F]=8'hFF;
    mem['h1F90]=8'hFF; mem['h1F91]=8'hFF; mem['h1F92]=8'hFF; mem['h1F93]=8'hFF;
    mem['h1F94]=8'hFF; mem['h1F95]=8'hFF; mem['h1F96]=8'hFF; mem['h1F97]=8'hFF;
    mem['h1F98]=8'hFF; mem['h1F99]=8'hFF; mem['h1F9A]=8'hFF; mem['h1F9B]=8'hFF;
    mem['h1F9C]=8'hFF; mem['h1F9D]=8'hFF; mem['h1F9E]=8'hFF; mem['h1F9F]=8'hFF;
    mem['h1FA0]=8'hFF; mem['h1FA1]=8'hFF; mem['h1FA2]=8'hFF; mem['h1FA3]=8'hFF;
    mem['h1FA4]=8'hFF; mem['h1FA5]=8'hFF; mem['h1FA6]=8'hFF; mem['h1FA7]=8'hFF;
    mem['h1FA8]=8'hFF; mem['h1FA9]=8'hFF; mem['h1FAA]=8'hFF; mem['h1FAB]=8'hFF;
    mem['h1FAC]=8'hFF; mem['h1FAD]=8'hFF; mem['h1FAE]=8'hFF; mem['h1FAF]=8'hFF;
    mem['h1FB0]=8'hFF; mem['h1FB1]=8'hFF; mem['h1FB2]=8'hFF; mem['h1FB3]=8'hFF;
    mem['h1FB4]=8'hFF; mem['h1FB5]=8'hFF; mem['h1FB6]=8'hFF; mem['h1FB7]=8'hFF;
    mem['h1FB8]=8'hFF; mem['h1FB9]=8'hFF; mem['h1FBA]=8'hFF; mem['h1FBB]=8'hFF;
    mem['h1FBC]=8'hFF; mem['h1FBD]=8'hFF; mem['h1FBE]=8'hFF; mem['h1FBF]=8'hFF;
    mem['h1FC0]=8'hFF; mem['h1FC1]=8'hFF; mem['h1FC2]=8'hFF; mem['h1FC3]=8'hFF;
    mem['h1FC4]=8'hFF; mem['h1FC5]=8'hFF; mem['h1FC6]=8'hFF; mem['h1FC7]=8'hFF;
    mem['h1FC8]=8'hFF; mem['h1FC9]=8'hFF; mem['h1FCA]=8'hFF; mem['h1FCB]=8'hFF;
    mem['h1FCC]=8'hFF; mem['h1FCD]=8'hFF; mem['h1FCE]=8'hFF; mem['h1FCF]=8'hFF;
    mem['h1FD0]=8'hFF; mem['h1FD1]=8'hFF; mem['h1FD2]=8'hFF; mem['h1FD3]=8'hFF;
    mem['h1FD4]=8'hFF; mem['h1FD5]=8'hFF; mem['h1FD6]=8'hFF; mem['h1FD7]=8'hFF;
    mem['h1FD8]=8'hFF; mem['h1FD9]=8'hFF; mem['h1FDA]=8'hFF; mem['h1FDB]=8'hFF;
    mem['h1FDC]=8'hFF; mem['h1FDD]=8'hFF; mem['h1FDE]=8'hFF; mem['h1FDF]=8'hFF;
    mem['h1FE0]=8'hFF; mem['h1FE1]=8'hFF; mem['h1FE2]=8'hFF; mem['h1FE3]=8'hFF;
    mem['h1FE4]=8'hFF; mem['h1FE5]=8'hFF; mem['h1FE6]=8'hFF; mem['h1FE7]=8'hFF;
    mem['h1FE8]=8'hFF; mem['h1FE9]=8'hFF; mem['h1FEA]=8'hFF; mem['h1FEB]=8'hFF;
    mem['h1FEC]=8'hFF; mem['h1FED]=8'hFF; mem['h1FEE]=8'hFF; mem['h1FEF]=8'hFF;
    mem['h1FF0]=8'hFF; mem['h1FF1]=8'hFF; mem['h1FF2]=8'hFF; mem['h1FF3]=8'hFF;
    mem['h1FF4]=8'hFF; mem['h1FF5]=8'hFF; mem['h1FF6]=8'hFF; mem['h1FF7]=8'hFF;
    mem['h1FF8]=8'hFF; mem['h1FF9]=8'hFF; mem['h1FFA]=8'hFF; mem['h1FFB]=8'hFF;
    mem['h1FFC]=8'hFF; mem['h1FFD]=8'hFF; mem['h1FFE]=8'hFF; mem['h1FFF]=8'hFF;
    mem['h2000]=8'hFF; mem['h2001]=8'hFF; mem['h2002]=8'hFF; mem['h2003]=8'hFF;
    mem['h2004]=8'hFF; mem['h2005]=8'hFF; mem['h2006]=8'hFF; mem['h2007]=8'hFF;
    mem['h2008]=8'hFF; mem['h2009]=8'hFF; mem['h200A]=8'hFF; mem['h200B]=8'hFF;
    mem['h200C]=8'hFF; mem['h200D]=8'hFF; mem['h200E]=8'hFF; mem['h200F]=8'hFF;
    mem['h2010]=8'hFF; mem['h2011]=8'hFF; mem['h2012]=8'hFF; mem['h2013]=8'hFF;
    mem['h2014]=8'hFF; mem['h2015]=8'hFF; mem['h2016]=8'hFF; mem['h2017]=8'hFF;
    mem['h2018]=8'hFF; mem['h2019]=8'hFF; mem['h201A]=8'hFF; mem['h201B]=8'hFF;
    mem['h201C]=8'hFF; mem['h201D]=8'hFF; mem['h201E]=8'hFF; mem['h201F]=8'hFF;
    mem['h2020]=8'hFF; mem['h2021]=8'hFF; mem['h2022]=8'hFF; mem['h2023]=8'hFF;
    mem['h2024]=8'hFF; mem['h2025]=8'hFF; mem['h2026]=8'hFF; mem['h2027]=8'hFF;
    mem['h2028]=8'hFF; mem['h2029]=8'hFF; mem['h202A]=8'hFF; mem['h202B]=8'hFF;
    mem['h202C]=8'hFF; mem['h202D]=8'hFF; mem['h202E]=8'hFF; mem['h202F]=8'hFF;
    mem['h2030]=8'hFF; mem['h2031]=8'hFF; mem['h2032]=8'hFF; mem['h2033]=8'hFF;
    mem['h2034]=8'hFF; mem['h2035]=8'hFF; mem['h2036]=8'hFF; mem['h2037]=8'hFF;
    mem['h2038]=8'hFF; mem['h2039]=8'hFF; mem['h203A]=8'hFF; mem['h203B]=8'hFF;
    mem['h203C]=8'hFF; mem['h203D]=8'hFF; mem['h203E]=8'hFF; mem['h203F]=8'hFF;
    mem['h2040]=8'hFF; mem['h2041]=8'hFF; mem['h2042]=8'hFF; mem['h2043]=8'hFF;
    mem['h2044]=8'hFF; mem['h2045]=8'hFF; mem['h2046]=8'hFF; mem['h2047]=8'hFF;
    mem['h2048]=8'hFF; mem['h2049]=8'hFF; mem['h204A]=8'hFF; mem['h204B]=8'hFF;
    mem['h204C]=8'hFF; mem['h204D]=8'hFF; mem['h204E]=8'hFF; mem['h204F]=8'hFF;
    mem['h2050]=8'hFF; mem['h2051]=8'hFF; mem['h2052]=8'hFF; mem['h2053]=8'hFF;
    mem['h2054]=8'hFF; mem['h2055]=8'hFF; mem['h2056]=8'hFF; mem['h2057]=8'hFF;
    mem['h2058]=8'hFF; mem['h2059]=8'hFF; mem['h205A]=8'hFF; mem['h205B]=8'hFF;
    mem['h205C]=8'hFF; mem['h205D]=8'hFF; mem['h205E]=8'hFF; mem['h205F]=8'hFF;
    mem['h2060]=8'hFF; mem['h2061]=8'hFF; mem['h2062]=8'hFF; mem['h2063]=8'hFF;
    mem['h2064]=8'hFF; mem['h2065]=8'hFF; mem['h2066]=8'hFF; mem['h2067]=8'hFF;
    mem['h2068]=8'hFF; mem['h2069]=8'hFF; mem['h206A]=8'hFF; mem['h206B]=8'hFF;
    mem['h206C]=8'hFF; mem['h206D]=8'hFF; mem['h206E]=8'hFF; mem['h206F]=8'hFF;
    mem['h2070]=8'hFF; mem['h2071]=8'hFF; mem['h2072]=8'hFF; mem['h2073]=8'hFF;
    mem['h2074]=8'hFF; mem['h2075]=8'hFF; mem['h2076]=8'hFF; mem['h2077]=8'hFF;
    mem['h2078]=8'hFF; mem['h2079]=8'hFF; mem['h207A]=8'hFF; mem['h207B]=8'hFF;
    mem['h207C]=8'hFF; mem['h207D]=8'hFF; mem['h207E]=8'hFF; mem['h207F]=8'hFF;
    mem['h2080]=8'hFF; mem['h2081]=8'hFF; mem['h2082]=8'hFF; mem['h2083]=8'hFF;
    mem['h2084]=8'hFF; mem['h2085]=8'hFF; mem['h2086]=8'hFF; mem['h2087]=8'hFF;
    mem['h2088]=8'hFF; mem['h2089]=8'hFF; mem['h208A]=8'hFF; mem['h208B]=8'hFF;
    mem['h208C]=8'hFF; mem['h208D]=8'hFF; mem['h208E]=8'hFF; mem['h208F]=8'hFF;
    mem['h2090]=8'hFF; mem['h2091]=8'hFF; mem['h2092]=8'hFF; mem['h2093]=8'hFF;
    mem['h2094]=8'hFF; mem['h2095]=8'hFF; mem['h2096]=8'hFF; mem['h2097]=8'hFF;
    mem['h2098]=8'hFF; mem['h2099]=8'hFF; mem['h209A]=8'hFF; mem['h209B]=8'hFF;
    mem['h209C]=8'hFF; mem['h209D]=8'hFF; mem['h209E]=8'hFF; mem['h209F]=8'hFF;
    mem['h20A0]=8'hFF; mem['h20A1]=8'hFF; mem['h20A2]=8'hFF; mem['h20A3]=8'hFF;
    mem['h20A4]=8'hFF; mem['h20A5]=8'hFF; mem['h20A6]=8'hFF; mem['h20A7]=8'hFF;
    mem['h20A8]=8'hFF; mem['h20A9]=8'hFF; mem['h20AA]=8'hFF; mem['h20AB]=8'hFF;
    mem['h20AC]=8'hFF; mem['h20AD]=8'hFF; mem['h20AE]=8'hFF; mem['h20AF]=8'hFF;
    mem['h20B0]=8'hFF; mem['h20B1]=8'hFF; mem['h20B2]=8'hFF; mem['h20B3]=8'hFF;
    mem['h20B4]=8'hFF; mem['h20B5]=8'hFF; mem['h20B6]=8'hFF; mem['h20B7]=8'hFF;
    mem['h20B8]=8'hFF; mem['h20B9]=8'hFF; mem['h20BA]=8'hFF; mem['h20BB]=8'hFF;
    mem['h20BC]=8'hFF; mem['h20BD]=8'hFF; mem['h20BE]=8'hFF; mem['h20BF]=8'hFF;
    mem['h20C0]=8'hFF; mem['h20C1]=8'hFF; mem['h20C2]=8'hFF; mem['h20C3]=8'hFF;
    mem['h20C4]=8'hFF; mem['h20C5]=8'hFF; mem['h20C6]=8'hFF; mem['h20C7]=8'hFF;
    mem['h20C8]=8'hFF; mem['h20C9]=8'hFF; mem['h20CA]=8'hFF; mem['h20CB]=8'hFF;
    mem['h20CC]=8'hFF; mem['h20CD]=8'hFF; mem['h20CE]=8'hFF; mem['h20CF]=8'hFF;
    mem['h20D0]=8'hFF; mem['h20D1]=8'hFF; mem['h20D2]=8'hFF; mem['h20D3]=8'hFF;
    mem['h20D4]=8'hFF; mem['h20D5]=8'hFF; mem['h20D6]=8'hFF; mem['h20D7]=8'hFF;
    mem['h20D8]=8'hFF; mem['h20D9]=8'hFF; mem['h20DA]=8'hFF; mem['h20DB]=8'hFF;
    mem['h20DC]=8'hFF; mem['h20DD]=8'hFF; mem['h20DE]=8'hFF; mem['h20DF]=8'hFF;
    mem['h20E0]=8'hFF; mem['h20E1]=8'hFF; mem['h20E2]=8'hFF; mem['h20E3]=8'hFF;
    mem['h20E4]=8'hFF; mem['h20E5]=8'hFF; mem['h20E6]=8'hFF; mem['h20E7]=8'hFF;
    mem['h20E8]=8'hFF; mem['h20E9]=8'hFF; mem['h20EA]=8'hFF; mem['h20EB]=8'hFF;
    mem['h20EC]=8'hFF; mem['h20ED]=8'hFF; mem['h20EE]=8'hFF; mem['h20EF]=8'hFF;
    mem['h20F0]=8'hFF; mem['h20F1]=8'hFF; mem['h20F2]=8'hFF; mem['h20F3]=8'hFF;
    mem['h20F4]=8'hFF; mem['h20F5]=8'hFF; mem['h20F6]=8'hFF; mem['h20F7]=8'hFF;
    mem['h20F8]=8'hFF; mem['h20F9]=8'hFF; mem['h20FA]=8'hFF; mem['h20FB]=8'hFF;
    mem['h20FC]=8'hFF; mem['h20FD]=8'hFF; mem['h20FE]=8'hFF; mem['h20FF]=8'hFF;
    mem['h2100]=8'hFF; mem['h2101]=8'hFF; mem['h2102]=8'hFF; mem['h2103]=8'hFF;
    mem['h2104]=8'hFF; mem['h2105]=8'hFF; mem['h2106]=8'hFF; mem['h2107]=8'hFF;
    mem['h2108]=8'hFF; mem['h2109]=8'hFF; mem['h210A]=8'hFF; mem['h210B]=8'hFF;
    mem['h210C]=8'hFF; mem['h210D]=8'hFF; mem['h210E]=8'hFF; mem['h210F]=8'hFF;
    mem['h2110]=8'hFF; mem['h2111]=8'hFF; mem['h2112]=8'hFF; mem['h2113]=8'hFF;
    mem['h2114]=8'hFF; mem['h2115]=8'hFF; mem['h2116]=8'hFF; mem['h2117]=8'hFF;
    mem['h2118]=8'hFF; mem['h2119]=8'hFF; mem['h211A]=8'hFF; mem['h211B]=8'hFF;
    mem['h211C]=8'hFF; mem['h211D]=8'hFF; mem['h211E]=8'hFF; mem['h211F]=8'hFF;
    mem['h2120]=8'hFF; mem['h2121]=8'hFF; mem['h2122]=8'hFF; mem['h2123]=8'hFF;
    mem['h2124]=8'hFF; mem['h2125]=8'hFF; mem['h2126]=8'hFF; mem['h2127]=8'hFF;
    mem['h2128]=8'hFF; mem['h2129]=8'hFF; mem['h212A]=8'hFF; mem['h212B]=8'hFF;
    mem['h212C]=8'hFF; mem['h212D]=8'hFF; mem['h212E]=8'hFF; mem['h212F]=8'hFF;
    mem['h2130]=8'hFF; mem['h2131]=8'hFF; mem['h2132]=8'hFF; mem['h2133]=8'hFF;
    mem['h2134]=8'hFF; mem['h2135]=8'hFF; mem['h2136]=8'hFF; mem['h2137]=8'hFF;
    mem['h2138]=8'hFF; mem['h2139]=8'hFF; mem['h213A]=8'hFF; mem['h213B]=8'hFF;
    mem['h213C]=8'hFF; mem['h213D]=8'hFF; mem['h213E]=8'hFF; mem['h213F]=8'hFF;
    mem['h2140]=8'hFF; mem['h2141]=8'hFF; mem['h2142]=8'hFF; mem['h2143]=8'hFF;
    mem['h2144]=8'hFF; mem['h2145]=8'hFF; mem['h2146]=8'hFF; mem['h2147]=8'hFF;
    mem['h2148]=8'hFF; mem['h2149]=8'hFF; mem['h214A]=8'hFF; mem['h214B]=8'hFF;
    mem['h214C]=8'hFF; mem['h214D]=8'hFF; mem['h214E]=8'hFF; mem['h214F]=8'hFF;
    mem['h2150]=8'hFF; mem['h2151]=8'hFF; mem['h2152]=8'hFF; mem['h2153]=8'hFF;
    mem['h2154]=8'hFF; mem['h2155]=8'hFF; mem['h2156]=8'hFF; mem['h2157]=8'hFF;
    mem['h2158]=8'hFF; mem['h2159]=8'hFF; mem['h215A]=8'hFF; mem['h215B]=8'hFF;
    mem['h215C]=8'hFF; mem['h215D]=8'hFF; mem['h215E]=8'hFF; mem['h215F]=8'hFF;
    mem['h2160]=8'hFF; mem['h2161]=8'hFF; mem['h2162]=8'hFF; mem['h2163]=8'hFF;
    mem['h2164]=8'hFF; mem['h2165]=8'hFF; mem['h2166]=8'hFF; mem['h2167]=8'hFF;
    mem['h2168]=8'hFF; mem['h2169]=8'hFF; mem['h216A]=8'hFF; mem['h216B]=8'hFF;
    mem['h216C]=8'hFF; mem['h216D]=8'hFF; mem['h216E]=8'hFF; mem['h216F]=8'hFF;
    mem['h2170]=8'hFF; mem['h2171]=8'hFF; mem['h2172]=8'hFF; mem['h2173]=8'hFF;
    mem['h2174]=8'hFF; mem['h2175]=8'hFF; mem['h2176]=8'hFF; mem['h2177]=8'hFF;
    mem['h2178]=8'hFF; mem['h2179]=8'hFF; mem['h217A]=8'hFF; mem['h217B]=8'hFF;
    mem['h217C]=8'hFF; mem['h217D]=8'hFF; mem['h217E]=8'hFF; mem['h217F]=8'hFF;
    mem['h2180]=8'hFF; mem['h2181]=8'hFF; mem['h2182]=8'hFF; mem['h2183]=8'hFF;
    mem['h2184]=8'hFF; mem['h2185]=8'hFF; mem['h2186]=8'hFF; mem['h2187]=8'hFF;
    mem['h2188]=8'hFF; mem['h2189]=8'hFF; mem['h218A]=8'hFF; mem['h218B]=8'hFF;
    mem['h218C]=8'hFF; mem['h218D]=8'hFF; mem['h218E]=8'hFF; mem['h218F]=8'hFF;
    mem['h2190]=8'hFF; mem['h2191]=8'hFF; mem['h2192]=8'hFF; mem['h2193]=8'hFF;
    mem['h2194]=8'hFF; mem['h2195]=8'hFF; mem['h2196]=8'hFF; mem['h2197]=8'hFF;
    mem['h2198]=8'hFF; mem['h2199]=8'hFF; mem['h219A]=8'hFF; mem['h219B]=8'hFF;
    mem['h219C]=8'hFF; mem['h219D]=8'hFF; mem['h219E]=8'hFF; mem['h219F]=8'hFF;
    mem['h21A0]=8'hFF; mem['h21A1]=8'hFF; mem['h21A2]=8'hFF; mem['h21A3]=8'hFF;
    mem['h21A4]=8'hFF; mem['h21A5]=8'hFF; mem['h21A6]=8'hFF; mem['h21A7]=8'hFF;
    mem['h21A8]=8'hFF; mem['h21A9]=8'hFF; mem['h21AA]=8'hFF; mem['h21AB]=8'hFF;
    mem['h21AC]=8'hFF; mem['h21AD]=8'hFF; mem['h21AE]=8'hFF; mem['h21AF]=8'hFF;
    mem['h21B0]=8'hFF; mem['h21B1]=8'hFF; mem['h21B2]=8'hFF; mem['h21B3]=8'hFF;
    mem['h21B4]=8'hFF; mem['h21B5]=8'hFF; mem['h21B6]=8'hFF; mem['h21B7]=8'hFF;
    mem['h21B8]=8'hFF; mem['h21B9]=8'hFF; mem['h21BA]=8'hFF; mem['h21BB]=8'hFF;
    mem['h21BC]=8'hFF; mem['h21BD]=8'hFF; mem['h21BE]=8'hFF; mem['h21BF]=8'hFF;
    mem['h21C0]=8'hFF; mem['h21C1]=8'hFF; mem['h21C2]=8'hFF; mem['h21C3]=8'hFF;
    mem['h21C4]=8'hFF; mem['h21C5]=8'hFF; mem['h21C6]=8'hFF; mem['h21C7]=8'hFF;
    mem['h21C8]=8'hFF; mem['h21C9]=8'hFF; mem['h21CA]=8'hFF; mem['h21CB]=8'hFF;
    mem['h21CC]=8'hFF; mem['h21CD]=8'hFF; mem['h21CE]=8'hFF; mem['h21CF]=8'hFF;
    mem['h21D0]=8'hFF; mem['h21D1]=8'hFF; mem['h21D2]=8'hFF; mem['h21D3]=8'hFF;
    mem['h21D4]=8'hFF; mem['h21D5]=8'hFF; mem['h21D6]=8'hFF; mem['h21D7]=8'hFF;
    mem['h21D8]=8'hFF; mem['h21D9]=8'hFF; mem['h21DA]=8'hFF; mem['h21DB]=8'hFF;
    mem['h21DC]=8'hFF; mem['h21DD]=8'hFF; mem['h21DE]=8'hFF; mem['h21DF]=8'hFF;
    mem['h21E0]=8'hFF; mem['h21E1]=8'hFF; mem['h21E2]=8'hFF; mem['h21E3]=8'hFF;
    mem['h21E4]=8'hFF; mem['h21E5]=8'hFF; mem['h21E6]=8'hFF; mem['h21E7]=8'hFF;
    mem['h21E8]=8'hFF; mem['h21E9]=8'hFF; mem['h21EA]=8'hFF; mem['h21EB]=8'hFF;
    mem['h21EC]=8'hFF; mem['h21ED]=8'hFF; mem['h21EE]=8'hFF; mem['h21EF]=8'hFF;
    mem['h21F0]=8'hFF; mem['h21F1]=8'hFF; mem['h21F2]=8'hFF; mem['h21F3]=8'hFF;
    mem['h21F4]=8'hFF; mem['h21F5]=8'hFF; mem['h21F6]=8'hFF; mem['h21F7]=8'hFF;
    mem['h21F8]=8'hFF; mem['h21F9]=8'hFF; mem['h21FA]=8'hFF; mem['h21FB]=8'hFF;
    mem['h21FC]=8'hFF; mem['h21FD]=8'hFF; mem['h21FE]=8'hFF; mem['h21FF]=8'hFF;
    mem['h2200]=8'hFF; mem['h2201]=8'hFF; mem['h2202]=8'hFF; mem['h2203]=8'hFF;
    mem['h2204]=8'hFF; mem['h2205]=8'hFF; mem['h2206]=8'hFF; mem['h2207]=8'hFF;
    mem['h2208]=8'hFF; mem['h2209]=8'hFF; mem['h220A]=8'hFF; mem['h220B]=8'hFF;
    mem['h220C]=8'hFF; mem['h220D]=8'hFF; mem['h220E]=8'hFF; mem['h220F]=8'hFF;
    mem['h2210]=8'hFF; mem['h2211]=8'hFF; mem['h2212]=8'hFF; mem['h2213]=8'hFF;
    mem['h2214]=8'hFF; mem['h2215]=8'hFF; mem['h2216]=8'hFF; mem['h2217]=8'hFF;
    mem['h2218]=8'hFF; mem['h2219]=8'hFF; mem['h221A]=8'hFF; mem['h221B]=8'hFF;
    mem['h221C]=8'hFF; mem['h221D]=8'hFF; mem['h221E]=8'hFF; mem['h221F]=8'hFF;
    mem['h2220]=8'hFF; mem['h2221]=8'hFF; mem['h2222]=8'hFF; mem['h2223]=8'hFF;
    mem['h2224]=8'hFF; mem['h2225]=8'hFF; mem['h2226]=8'hFF; mem['h2227]=8'hFF;
    mem['h2228]=8'hFF; mem['h2229]=8'hFF; mem['h222A]=8'hFF; mem['h222B]=8'hFF;
    mem['h222C]=8'hFF; mem['h222D]=8'hFF; mem['h222E]=8'hFF; mem['h222F]=8'hFF;
    mem['h2230]=8'hFF; mem['h2231]=8'hFF; mem['h2232]=8'hFF; mem['h2233]=8'hFF;
    mem['h2234]=8'hFF; mem['h2235]=8'hFF; mem['h2236]=8'hFF; mem['h2237]=8'hFF;
    mem['h2238]=8'hFF; mem['h2239]=8'hFF; mem['h223A]=8'hFF; mem['h223B]=8'hFF;
    mem['h223C]=8'hFF; mem['h223D]=8'hFF; mem['h223E]=8'hFF; mem['h223F]=8'hFF;
    mem['h2240]=8'hFF; mem['h2241]=8'hFF; mem['h2242]=8'hFF; mem['h2243]=8'hFF;
    mem['h2244]=8'hFF; mem['h2245]=8'hFF; mem['h2246]=8'hFF; mem['h2247]=8'hFF;
    mem['h2248]=8'hFF; mem['h2249]=8'hFF; mem['h224A]=8'hFF; mem['h224B]=8'hFF;
    mem['h224C]=8'hFF; mem['h224D]=8'hFF; mem['h224E]=8'hFF; mem['h224F]=8'hFF;
    mem['h2250]=8'hFF; mem['h2251]=8'hFF; mem['h2252]=8'hFF; mem['h2253]=8'hFF;
    mem['h2254]=8'hFF; mem['h2255]=8'hFF; mem['h2256]=8'hFF; mem['h2257]=8'hFF;
    mem['h2258]=8'hFF; mem['h2259]=8'hFF; mem['h225A]=8'hFF; mem['h225B]=8'hFF;
    mem['h225C]=8'hFF; mem['h225D]=8'hFF; mem['h225E]=8'hFF; mem['h225F]=8'hFF;
    mem['h2260]=8'hFF; mem['h2261]=8'hFF; mem['h2262]=8'hFF; mem['h2263]=8'hFF;
    mem['h2264]=8'hFF; mem['h2265]=8'hFF; mem['h2266]=8'hFF; mem['h2267]=8'hFF;
    mem['h2268]=8'hFF; mem['h2269]=8'hFF; mem['h226A]=8'hFF; mem['h226B]=8'hFF;
    mem['h226C]=8'hFF; mem['h226D]=8'hFF; mem['h226E]=8'hFF; mem['h226F]=8'hFF;
    mem['h2270]=8'hFF; mem['h2271]=8'hFF; mem['h2272]=8'hFF; mem['h2273]=8'hFF;
    mem['h2274]=8'hFF; mem['h2275]=8'hFF; mem['h2276]=8'hFF; mem['h2277]=8'hFF;
    mem['h2278]=8'hFF; mem['h2279]=8'hFF; mem['h227A]=8'hFF; mem['h227B]=8'hFF;
    mem['h227C]=8'hFF; mem['h227D]=8'hFF; mem['h227E]=8'hFF; mem['h227F]=8'hFF;
    mem['h2280]=8'hFF; mem['h2281]=8'hFF; mem['h2282]=8'hFF; mem['h2283]=8'hFF;
    mem['h2284]=8'hFF; mem['h2285]=8'hFF; mem['h2286]=8'hFF; mem['h2287]=8'hFF;
    mem['h2288]=8'hFF; mem['h2289]=8'hFF; mem['h228A]=8'hFF; mem['h228B]=8'hFF;
    mem['h228C]=8'hFF; mem['h228D]=8'hFF; mem['h228E]=8'hFF; mem['h228F]=8'hFF;
    mem['h2290]=8'hFF; mem['h2291]=8'hFF; mem['h2292]=8'hFF; mem['h2293]=8'hFF;
    mem['h2294]=8'hFF; mem['h2295]=8'hFF; mem['h2296]=8'hFF; mem['h2297]=8'hFF;
    mem['h2298]=8'hFF; mem['h2299]=8'hFF; mem['h229A]=8'hFF; mem['h229B]=8'hFF;
    mem['h229C]=8'hFF; mem['h229D]=8'hFF; mem['h229E]=8'hFF; mem['h229F]=8'hFF;
    mem['h22A0]=8'hFF; mem['h22A1]=8'hFF; mem['h22A2]=8'hFF; mem['h22A3]=8'hFF;
    mem['h22A4]=8'hFF; mem['h22A5]=8'hFF; mem['h22A6]=8'hFF; mem['h22A7]=8'hFF;
    mem['h22A8]=8'hFF; mem['h22A9]=8'hFF; mem['h22AA]=8'hFF; mem['h22AB]=8'hFF;
    mem['h22AC]=8'hFF; mem['h22AD]=8'hFF; mem['h22AE]=8'hFF; mem['h22AF]=8'hFF;
    mem['h22B0]=8'hFF; mem['h22B1]=8'hFF; mem['h22B2]=8'hFF; mem['h22B3]=8'hFF;
    mem['h22B4]=8'hFF; mem['h22B5]=8'hFF; mem['h22B6]=8'hFF; mem['h22B7]=8'hFF;
    mem['h22B8]=8'hFF; mem['h22B9]=8'hFF; mem['h22BA]=8'hFF; mem['h22BB]=8'hFF;
    mem['h22BC]=8'hFF; mem['h22BD]=8'hFF; mem['h22BE]=8'hFF; mem['h22BF]=8'hFF;
    mem['h22C0]=8'hFF; mem['h22C1]=8'hFF; mem['h22C2]=8'hFF; mem['h22C3]=8'hFF;
    mem['h22C4]=8'hFF; mem['h22C5]=8'hFF; mem['h22C6]=8'hFF; mem['h22C7]=8'hFF;
    mem['h22C8]=8'hFF; mem['h22C9]=8'hFF; mem['h22CA]=8'hFF; mem['h22CB]=8'hFF;
    mem['h22CC]=8'hFF; mem['h22CD]=8'hFF; mem['h22CE]=8'hFF; mem['h22CF]=8'hFF;
    mem['h22D0]=8'hFF; mem['h22D1]=8'hFF; mem['h22D2]=8'hFF; mem['h22D3]=8'hFF;
    mem['h22D4]=8'hFF; mem['h22D5]=8'hFF; mem['h22D6]=8'hFF; mem['h22D7]=8'hFF;
    mem['h22D8]=8'hFF; mem['h22D9]=8'hFF; mem['h22DA]=8'hFF; mem['h22DB]=8'hFF;
    mem['h22DC]=8'hFF; mem['h22DD]=8'hFF; mem['h22DE]=8'hFF; mem['h22DF]=8'hFF;
    mem['h22E0]=8'hFF; mem['h22E1]=8'hFF; mem['h22E2]=8'hFF; mem['h22E3]=8'hFF;
    mem['h22E4]=8'hFF; mem['h22E5]=8'hFF; mem['h22E6]=8'hFF; mem['h22E7]=8'hFF;
    mem['h22E8]=8'hFF; mem['h22E9]=8'hFF; mem['h22EA]=8'hFF; mem['h22EB]=8'hFF;
    mem['h22EC]=8'hFF; mem['h22ED]=8'hFF; mem['h22EE]=8'hFF; mem['h22EF]=8'hFF;
    mem['h22F0]=8'hFF; mem['h22F1]=8'hFF; mem['h22F2]=8'hFF; mem['h22F3]=8'hFF;
    mem['h22F4]=8'hFF; mem['h22F5]=8'hFF; mem['h22F6]=8'hFF; mem['h22F7]=8'hFF;
    mem['h22F8]=8'hFF; mem['h22F9]=8'hFF; mem['h22FA]=8'hFF; mem['h22FB]=8'hFF;
    mem['h22FC]=8'hFF; mem['h22FD]=8'hFF; mem['h22FE]=8'hFF; mem['h22FF]=8'hFF;
    mem['h2300]=8'hFF; mem['h2301]=8'hFF; mem['h2302]=8'hFF; mem['h2303]=8'hFF;
    mem['h2304]=8'hFF; mem['h2305]=8'hFF; mem['h2306]=8'hFF; mem['h2307]=8'hFF;
    mem['h2308]=8'hFF; mem['h2309]=8'hFF; mem['h230A]=8'hFF; mem['h230B]=8'hFF;
    mem['h230C]=8'hFF; mem['h230D]=8'hFF; mem['h230E]=8'hFF; mem['h230F]=8'hFF;
    mem['h2310]=8'hFF; mem['h2311]=8'hFF; mem['h2312]=8'hFF; mem['h2313]=8'hFF;
    mem['h2314]=8'hFF; mem['h2315]=8'hFF; mem['h2316]=8'hFF; mem['h2317]=8'hFF;
    mem['h2318]=8'hFF; mem['h2319]=8'hFF; mem['h231A]=8'hFF; mem['h231B]=8'hFF;
    mem['h231C]=8'hFF; mem['h231D]=8'hFF; mem['h231E]=8'hFF; mem['h231F]=8'hFF;
    mem['h2320]=8'hFF; mem['h2321]=8'hFF; mem['h2322]=8'hFF; mem['h2323]=8'hFF;
    mem['h2324]=8'hFF; mem['h2325]=8'hFF; mem['h2326]=8'hFF; mem['h2327]=8'hFF;
    mem['h2328]=8'hFF; mem['h2329]=8'hFF; mem['h232A]=8'hFF; mem['h232B]=8'hFF;
    mem['h232C]=8'hFF; mem['h232D]=8'hFF; mem['h232E]=8'hFF; mem['h232F]=8'hFF;
    mem['h2330]=8'hFF; mem['h2331]=8'hFF; mem['h2332]=8'hFF; mem['h2333]=8'hFF;
    mem['h2334]=8'hFF; mem['h2335]=8'hFF; mem['h2336]=8'hFF; mem['h2337]=8'hFF;
    mem['h2338]=8'hFF; mem['h2339]=8'hFF; mem['h233A]=8'hFF; mem['h233B]=8'hFF;
    mem['h233C]=8'hFF; mem['h233D]=8'hFF; mem['h233E]=8'hFF; mem['h233F]=8'hFF;
    mem['h2340]=8'hFF; mem['h2341]=8'hFF; mem['h2342]=8'hFF; mem['h2343]=8'hFF;
    mem['h2344]=8'hFF; mem['h2345]=8'hFF; mem['h2346]=8'hFF; mem['h2347]=8'hFF;
    mem['h2348]=8'hFF; mem['h2349]=8'hFF; mem['h234A]=8'hFF; mem['h234B]=8'hFF;
    mem['h234C]=8'hFF; mem['h234D]=8'hFF; mem['h234E]=8'hFF; mem['h234F]=8'hFF;
    mem['h2350]=8'hFF; mem['h2351]=8'hFF; mem['h2352]=8'hFF; mem['h2353]=8'hFF;
    mem['h2354]=8'hFF; mem['h2355]=8'hFF; mem['h2356]=8'hFF; mem['h2357]=8'hFF;
    mem['h2358]=8'hFF; mem['h2359]=8'hFF; mem['h235A]=8'hFF; mem['h235B]=8'hFF;
    mem['h235C]=8'hFF; mem['h235D]=8'hFF; mem['h235E]=8'hFF; mem['h235F]=8'hFF;
    mem['h2360]=8'hFF; mem['h2361]=8'hFF; mem['h2362]=8'hFF; mem['h2363]=8'hFF;
    mem['h2364]=8'hFF; mem['h2365]=8'hFF; mem['h2366]=8'hFF; mem['h2367]=8'hFF;
    mem['h2368]=8'hFF; mem['h2369]=8'hFF; mem['h236A]=8'hFF; mem['h236B]=8'hFF;
    mem['h236C]=8'hFF; mem['h236D]=8'hFF; mem['h236E]=8'hFF; mem['h236F]=8'hFF;
    mem['h2370]=8'hFF; mem['h2371]=8'hFF; mem['h2372]=8'hFF; mem['h2373]=8'hFF;
    mem['h2374]=8'hFF; mem['h2375]=8'hFF; mem['h2376]=8'hFF; mem['h2377]=8'hFF;
    mem['h2378]=8'hFF; mem['h2379]=8'hFF; mem['h237A]=8'hFF; mem['h237B]=8'hFF;
    mem['h237C]=8'hFF; mem['h237D]=8'hFF; mem['h237E]=8'hFF; mem['h237F]=8'hFF;
    mem['h2380]=8'hFF; mem['h2381]=8'hFF; mem['h2382]=8'hFF; mem['h2383]=8'hFF;
    mem['h2384]=8'hFF; mem['h2385]=8'hFF; mem['h2386]=8'hFF; mem['h2387]=8'hFF;
    mem['h2388]=8'hFF; mem['h2389]=8'hFF; mem['h238A]=8'hFF; mem['h238B]=8'hFF;
    mem['h238C]=8'hFF; mem['h238D]=8'hFF; mem['h238E]=8'hFF; mem['h238F]=8'hFF;
    mem['h2390]=8'hFF; mem['h2391]=8'hFF; mem['h2392]=8'hFF; mem['h2393]=8'hFF;
    mem['h2394]=8'hFF; mem['h2395]=8'hFF; mem['h2396]=8'hFF; mem['h2397]=8'hFF;
    mem['h2398]=8'hFF; mem['h2399]=8'hFF; mem['h239A]=8'hFF; mem['h239B]=8'hFF;
    mem['h239C]=8'hFF; mem['h239D]=8'hFF; mem['h239E]=8'hFF; mem['h239F]=8'hFF;
    mem['h23A0]=8'hFF; mem['h23A1]=8'hFF; mem['h23A2]=8'hFF; mem['h23A3]=8'hFF;
    mem['h23A4]=8'hFF; mem['h23A5]=8'hFF; mem['h23A6]=8'hFF; mem['h23A7]=8'hFF;
    mem['h23A8]=8'hFF; mem['h23A9]=8'hFF; mem['h23AA]=8'hFF; mem['h23AB]=8'hFF;
    mem['h23AC]=8'hFF; mem['h23AD]=8'hFF; mem['h23AE]=8'hFF; mem['h23AF]=8'hFF;
    mem['h23B0]=8'hFF; mem['h23B1]=8'hFF; mem['h23B2]=8'hFF; mem['h23B3]=8'hFF;
    mem['h23B4]=8'hFF; mem['h23B5]=8'hFF; mem['h23B6]=8'hFF; mem['h23B7]=8'hFF;
    mem['h23B8]=8'hFF; mem['h23B9]=8'hFF; mem['h23BA]=8'hFF; mem['h23BB]=8'hFF;
    mem['h23BC]=8'hFF; mem['h23BD]=8'hFF; mem['h23BE]=8'hFF; mem['h23BF]=8'hFF;
    mem['h23C0]=8'hFF; mem['h23C1]=8'hFF; mem['h23C2]=8'hFF; mem['h23C3]=8'hFF;
    mem['h23C4]=8'hFF; mem['h23C5]=8'hFF; mem['h23C6]=8'hFF; mem['h23C7]=8'hFF;
    mem['h23C8]=8'hFF; mem['h23C9]=8'hFF; mem['h23CA]=8'hFF; mem['h23CB]=8'hFF;
    mem['h23CC]=8'hFF; mem['h23CD]=8'hFF; mem['h23CE]=8'hFF; mem['h23CF]=8'hFF;
    mem['h23D0]=8'hFF; mem['h23D1]=8'hFF; mem['h23D2]=8'hFF; mem['h23D3]=8'hFF;
    mem['h23D4]=8'hFF; mem['h23D5]=8'hFF; mem['h23D6]=8'hFF; mem['h23D7]=8'hFF;
    mem['h23D8]=8'hFF; mem['h23D9]=8'hFF; mem['h23DA]=8'hFF; mem['h23DB]=8'hFF;
    mem['h23DC]=8'hFF; mem['h23DD]=8'hFF; mem['h23DE]=8'hFF; mem['h23DF]=8'hFF;
    mem['h23E0]=8'hFF; mem['h23E1]=8'hFF; mem['h23E2]=8'hFF; mem['h23E3]=8'hFF;
    mem['h23E4]=8'hFF; mem['h23E5]=8'hFF; mem['h23E6]=8'hFF; mem['h23E7]=8'hFF;
    mem['h23E8]=8'hFF; mem['h23E9]=8'hFF; mem['h23EA]=8'hFF; mem['h23EB]=8'hFF;
    mem['h23EC]=8'hFF; mem['h23ED]=8'hFF; mem['h23EE]=8'hFF; mem['h23EF]=8'hFF;
    mem['h23F0]=8'hFF; mem['h23F1]=8'hFF; mem['h23F2]=8'hFF; mem['h23F3]=8'hFF;
    mem['h23F4]=8'hFF; mem['h23F5]=8'hFF; mem['h23F6]=8'hFF; mem['h23F7]=8'hFF;
    mem['h23F8]=8'hFF; mem['h23F9]=8'hFF; mem['h23FA]=8'hFF; mem['h23FB]=8'hFF;
    mem['h23FC]=8'hFF; mem['h23FD]=8'hFF; mem['h23FE]=8'hFF; mem['h23FF]=8'hFF;
    mem['h2400]=8'hFF; mem['h2401]=8'hFF; mem['h2402]=8'hFF; mem['h2403]=8'hFF;
    mem['h2404]=8'hFF; mem['h2405]=8'hFF; mem['h2406]=8'hFF; mem['h2407]=8'hFF;
    mem['h2408]=8'hFF; mem['h2409]=8'hFF; mem['h240A]=8'hFF; mem['h240B]=8'hFF;
    mem['h240C]=8'hFF; mem['h240D]=8'hFF; mem['h240E]=8'hFF; mem['h240F]=8'hFF;
    mem['h2410]=8'hFF; mem['h2411]=8'hFF; mem['h2412]=8'hFF; mem['h2413]=8'hFF;
    mem['h2414]=8'hFF; mem['h2415]=8'hFF; mem['h2416]=8'hFF; mem['h2417]=8'hFF;
    mem['h2418]=8'hFF; mem['h2419]=8'hFF; mem['h241A]=8'hFF; mem['h241B]=8'hFF;
    mem['h241C]=8'hFF; mem['h241D]=8'hFF; mem['h241E]=8'hFF; mem['h241F]=8'hFF;
    mem['h2420]=8'hFF; mem['h2421]=8'hFF; mem['h2422]=8'hFF; mem['h2423]=8'hFF;
    mem['h2424]=8'hFF; mem['h2425]=8'hFF; mem['h2426]=8'hFF; mem['h2427]=8'hFF;
    mem['h2428]=8'hFF; mem['h2429]=8'hFF; mem['h242A]=8'hFF; mem['h242B]=8'hFF;
    mem['h242C]=8'hFF; mem['h242D]=8'hFF; mem['h242E]=8'hFF; mem['h242F]=8'hFF;
    mem['h2430]=8'hFF; mem['h2431]=8'hFF; mem['h2432]=8'hFF; mem['h2433]=8'hFF;
    mem['h2434]=8'hFF; mem['h2435]=8'hFF; mem['h2436]=8'hFF; mem['h2437]=8'hFF;
    mem['h2438]=8'hFF; mem['h2439]=8'hFF; mem['h243A]=8'hFF; mem['h243B]=8'hFF;
    mem['h243C]=8'hFF; mem['h243D]=8'hFF; mem['h243E]=8'hFF; mem['h243F]=8'hFF;
    mem['h2440]=8'hFF; mem['h2441]=8'hFF; mem['h2442]=8'hFF; mem['h2443]=8'hFF;
    mem['h2444]=8'hFF; mem['h2445]=8'hFF; mem['h2446]=8'hFF; mem['h2447]=8'hFF;
    mem['h2448]=8'hFF; mem['h2449]=8'hFF; mem['h244A]=8'hFF; mem['h244B]=8'hFF;
    mem['h244C]=8'hFF; mem['h244D]=8'hFF; mem['h244E]=8'hFF; mem['h244F]=8'hFF;
    mem['h2450]=8'hFF; mem['h2451]=8'hFF; mem['h2452]=8'hFF; mem['h2453]=8'hFF;
    mem['h2454]=8'hFF; mem['h2455]=8'hFF; mem['h2456]=8'hFF; mem['h2457]=8'hFF;
    mem['h2458]=8'hFF; mem['h2459]=8'hFF; mem['h245A]=8'hFF; mem['h245B]=8'hFF;
    mem['h245C]=8'hFF; mem['h245D]=8'hFF; mem['h245E]=8'hFF; mem['h245F]=8'hFF;
    mem['h2460]=8'hFF; mem['h2461]=8'hFF; mem['h2462]=8'hFF; mem['h2463]=8'hFF;
    mem['h2464]=8'hFF; mem['h2465]=8'hFF; mem['h2466]=8'hFF; mem['h2467]=8'hFF;
    mem['h2468]=8'hFF; mem['h2469]=8'hFF; mem['h246A]=8'hFF; mem['h246B]=8'hFF;
    mem['h246C]=8'hFF; mem['h246D]=8'hFF; mem['h246E]=8'hFF; mem['h246F]=8'hFF;
    mem['h2470]=8'hFF; mem['h2471]=8'hFF; mem['h2472]=8'hFF; mem['h2473]=8'hFF;
    mem['h2474]=8'hFF; mem['h2475]=8'hFF; mem['h2476]=8'hFF; mem['h2477]=8'hFF;
    mem['h2478]=8'hFF; mem['h2479]=8'hFF; mem['h247A]=8'hFF; mem['h247B]=8'hFF;
    mem['h247C]=8'hFF; mem['h247D]=8'hFF; mem['h247E]=8'hFF; mem['h247F]=8'hFF;
    mem['h2480]=8'hFF; mem['h2481]=8'hFF; mem['h2482]=8'hFF; mem['h2483]=8'hFF;
    mem['h2484]=8'hFF; mem['h2485]=8'hFF; mem['h2486]=8'hFF; mem['h2487]=8'hFF;
    mem['h2488]=8'hFF; mem['h2489]=8'hFF; mem['h248A]=8'hFF; mem['h248B]=8'hFF;
    mem['h248C]=8'hFF; mem['h248D]=8'hFF; mem['h248E]=8'hFF; mem['h248F]=8'hFF;
    mem['h2490]=8'hFF; mem['h2491]=8'hFF; mem['h2492]=8'hFF; mem['h2493]=8'hFF;
    mem['h2494]=8'hFF; mem['h2495]=8'hFF; mem['h2496]=8'hFF; mem['h2497]=8'hFF;
    mem['h2498]=8'hFF; mem['h2499]=8'hFF; mem['h249A]=8'hFF; mem['h249B]=8'hFF;
    mem['h249C]=8'hFF; mem['h249D]=8'hFF; mem['h249E]=8'hFF; mem['h249F]=8'hFF;
    mem['h24A0]=8'hFF; mem['h24A1]=8'hFF; mem['h24A2]=8'hFF; mem['h24A3]=8'hFF;
    mem['h24A4]=8'hFF; mem['h24A5]=8'hFF; mem['h24A6]=8'hFF; mem['h24A7]=8'hFF;
    mem['h24A8]=8'hFF; mem['h24A9]=8'hFF; mem['h24AA]=8'hFF; mem['h24AB]=8'hFF;
    mem['h24AC]=8'hFF; mem['h24AD]=8'hFF; mem['h24AE]=8'hFF; mem['h24AF]=8'hFF;
    mem['h24B0]=8'hFF; mem['h24B1]=8'hFF; mem['h24B2]=8'hFF; mem['h24B3]=8'hFF;
    mem['h24B4]=8'hFF; mem['h24B5]=8'hFF; mem['h24B6]=8'hFF; mem['h24B7]=8'hFF;
    mem['h24B8]=8'hFF; mem['h24B9]=8'hFF; mem['h24BA]=8'hFF; mem['h24BB]=8'hFF;
    mem['h24BC]=8'hFF; mem['h24BD]=8'hFF; mem['h24BE]=8'hFF; mem['h24BF]=8'hFF;
    mem['h24C0]=8'hFF; mem['h24C1]=8'hFF; mem['h24C2]=8'hFF; mem['h24C3]=8'hFF;
    mem['h24C4]=8'hFF; mem['h24C5]=8'hFF; mem['h24C6]=8'hFF; mem['h24C7]=8'hFF;
    mem['h24C8]=8'hFF; mem['h24C9]=8'hFF; mem['h24CA]=8'hFF; mem['h24CB]=8'hFF;
    mem['h24CC]=8'hFF; mem['h24CD]=8'hFF; mem['h24CE]=8'hFF; mem['h24CF]=8'hFF;
    mem['h24D0]=8'hFF; mem['h24D1]=8'hFF; mem['h24D2]=8'hFF; mem['h24D3]=8'hFF;
    mem['h24D4]=8'hFF; mem['h24D5]=8'hFF; mem['h24D6]=8'hFF; mem['h24D7]=8'hFF;
    mem['h24D8]=8'hFF; mem['h24D9]=8'hFF; mem['h24DA]=8'hFF; mem['h24DB]=8'hFF;
    mem['h24DC]=8'hFF; mem['h24DD]=8'hFF; mem['h24DE]=8'hFF; mem['h24DF]=8'hFF;
    mem['h24E0]=8'hFF; mem['h24E1]=8'hFF; mem['h24E2]=8'hFF; mem['h24E3]=8'hFF;
    mem['h24E4]=8'hFF; mem['h24E5]=8'hFF; mem['h24E6]=8'hFF; mem['h24E7]=8'hFF;
    mem['h24E8]=8'hFF; mem['h24E9]=8'hFF; mem['h24EA]=8'hFF; mem['h24EB]=8'hFF;
    mem['h24EC]=8'hFF; mem['h24ED]=8'hFF; mem['h24EE]=8'hFF; mem['h24EF]=8'hFF;
    mem['h24F0]=8'hFF; mem['h24F1]=8'hFF; mem['h24F2]=8'hFF; mem['h24F3]=8'hFF;
    mem['h24F4]=8'hFF; mem['h24F5]=8'hFF; mem['h24F6]=8'hFF; mem['h24F7]=8'hFF;
    mem['h24F8]=8'hFF; mem['h24F9]=8'hFF; mem['h24FA]=8'hFF; mem['h24FB]=8'hFF;
    mem['h24FC]=8'hFF; mem['h24FD]=8'hFF; mem['h24FE]=8'hFF; mem['h24FF]=8'hFF;
    mem['h2500]=8'hFF; mem['h2501]=8'hFF; mem['h2502]=8'hFF; mem['h2503]=8'hFF;
    mem['h2504]=8'hFF; mem['h2505]=8'hFF; mem['h2506]=8'hFF; mem['h2507]=8'hFF;
    mem['h2508]=8'hFF; mem['h2509]=8'hFF; mem['h250A]=8'hFF; mem['h250B]=8'hFF;
    mem['h250C]=8'hFF; mem['h250D]=8'hFF; mem['h250E]=8'hFF; mem['h250F]=8'hFF;
    mem['h2510]=8'hFF; mem['h2511]=8'hFF; mem['h2512]=8'hFF; mem['h2513]=8'hFF;
    mem['h2514]=8'hFF; mem['h2515]=8'hFF; mem['h2516]=8'hFF; mem['h2517]=8'hFF;
    mem['h2518]=8'hFF; mem['h2519]=8'hFF; mem['h251A]=8'hFF; mem['h251B]=8'hFF;
    mem['h251C]=8'hFF; mem['h251D]=8'hFF; mem['h251E]=8'hFF; mem['h251F]=8'hFF;
    mem['h2520]=8'hFF; mem['h2521]=8'hFF; mem['h2522]=8'hFF; mem['h2523]=8'hFF;
    mem['h2524]=8'hFF; mem['h2525]=8'hFF; mem['h2526]=8'hFF; mem['h2527]=8'hFF;
    mem['h2528]=8'hFF; mem['h2529]=8'hFF; mem['h252A]=8'hFF; mem['h252B]=8'hFF;
    mem['h252C]=8'hFF; mem['h252D]=8'hFF; mem['h252E]=8'hFF; mem['h252F]=8'hFF;
    mem['h2530]=8'hFF; mem['h2531]=8'hFF; mem['h2532]=8'hFF; mem['h2533]=8'hFF;
    mem['h2534]=8'hFF; mem['h2535]=8'hFF; mem['h2536]=8'hFF; mem['h2537]=8'hFF;
    mem['h2538]=8'hFF; mem['h2539]=8'hFF; mem['h253A]=8'hFF; mem['h253B]=8'hFF;
    mem['h253C]=8'hFF; mem['h253D]=8'hFF; mem['h253E]=8'hFF; mem['h253F]=8'hFF;
    mem['h2540]=8'hFF; mem['h2541]=8'hFF; mem['h2542]=8'hFF; mem['h2543]=8'hFF;
    mem['h2544]=8'hFF; mem['h2545]=8'hFF; mem['h2546]=8'hFF; mem['h2547]=8'hFF;
    mem['h2548]=8'hFF; mem['h2549]=8'hFF; mem['h254A]=8'hFF; mem['h254B]=8'hFF;
    mem['h254C]=8'hFF; mem['h254D]=8'hFF; mem['h254E]=8'hFF; mem['h254F]=8'hFF;
    mem['h2550]=8'hFF; mem['h2551]=8'hFF; mem['h2552]=8'hFF; mem['h2553]=8'hFF;
    mem['h2554]=8'hFF; mem['h2555]=8'hFF; mem['h2556]=8'hFF; mem['h2557]=8'hFF;
    mem['h2558]=8'hFF; mem['h2559]=8'hFF; mem['h255A]=8'hFF; mem['h255B]=8'hFF;
    mem['h255C]=8'hFF; mem['h255D]=8'hFF; mem['h255E]=8'hFF; mem['h255F]=8'hFF;
    mem['h2560]=8'hFF; mem['h2561]=8'hFF; mem['h2562]=8'hFF; mem['h2563]=8'hFF;
    mem['h2564]=8'hFF; mem['h2565]=8'hFF; mem['h2566]=8'hFF; mem['h2567]=8'hFF;
    mem['h2568]=8'hFF; mem['h2569]=8'hFF; mem['h256A]=8'hFF; mem['h256B]=8'hFF;
    mem['h256C]=8'hFF; mem['h256D]=8'hFF; mem['h256E]=8'hFF; mem['h256F]=8'hFF;
    mem['h2570]=8'hFF; mem['h2571]=8'hFF; mem['h2572]=8'hFF; mem['h2573]=8'hFF;
    mem['h2574]=8'hFF; mem['h2575]=8'hFF; mem['h2576]=8'hFF; mem['h2577]=8'hFF;
    mem['h2578]=8'hFF; mem['h2579]=8'hFF; mem['h257A]=8'hFF; mem['h257B]=8'hFF;
    mem['h257C]=8'hFF; mem['h257D]=8'hFF; mem['h257E]=8'hFF; mem['h257F]=8'hFF;
    mem['h2580]=8'hFF; mem['h2581]=8'hFF; mem['h2582]=8'hFF; mem['h2583]=8'hFF;
    mem['h2584]=8'hFF; mem['h2585]=8'hFF; mem['h2586]=8'hFF; mem['h2587]=8'hFF;
    mem['h2588]=8'hFF; mem['h2589]=8'hFF; mem['h258A]=8'hFF; mem['h258B]=8'hFF;
    mem['h258C]=8'hFF; mem['h258D]=8'hFF; mem['h258E]=8'hFF; mem['h258F]=8'hFF;
    mem['h2590]=8'hFF; mem['h2591]=8'hFF; mem['h2592]=8'hFF; mem['h2593]=8'hFF;
    mem['h2594]=8'hFF; mem['h2595]=8'hFF; mem['h2596]=8'hFF; mem['h2597]=8'hFF;
    mem['h2598]=8'hFF; mem['h2599]=8'hFF; mem['h259A]=8'hFF; mem['h259B]=8'hFF;
    mem['h259C]=8'hFF; mem['h259D]=8'hFF; mem['h259E]=8'hFF; mem['h259F]=8'hFF;
    mem['h25A0]=8'hFF; mem['h25A1]=8'hFF; mem['h25A2]=8'hFF; mem['h25A3]=8'hFF;
    mem['h25A4]=8'hFF; mem['h25A5]=8'hFF; mem['h25A6]=8'hFF; mem['h25A7]=8'hFF;
    mem['h25A8]=8'hFF; mem['h25A9]=8'hFF; mem['h25AA]=8'hFF; mem['h25AB]=8'hFF;
    mem['h25AC]=8'hFF; mem['h25AD]=8'hFF; mem['h25AE]=8'hFF; mem['h25AF]=8'hFF;
    mem['h25B0]=8'hFF; mem['h25B1]=8'hFF; mem['h25B2]=8'hFF; mem['h25B3]=8'hFF;
    mem['h25B4]=8'hFF; mem['h25B5]=8'hFF; mem['h25B6]=8'hFF; mem['h25B7]=8'hFF;
    mem['h25B8]=8'hFF; mem['h25B9]=8'hFF; mem['h25BA]=8'hFF; mem['h25BB]=8'hFF;
    mem['h25BC]=8'hFF; mem['h25BD]=8'hFF; mem['h25BE]=8'hFF; mem['h25BF]=8'hFF;
    mem['h25C0]=8'hFF; mem['h25C1]=8'hFF; mem['h25C2]=8'hFF; mem['h25C3]=8'hFF;
    mem['h25C4]=8'hFF; mem['h25C5]=8'hFF; mem['h25C6]=8'hFF; mem['h25C7]=8'hFF;
    mem['h25C8]=8'hFF; mem['h25C9]=8'hFF; mem['h25CA]=8'hFF; mem['h25CB]=8'hFF;
    mem['h25CC]=8'hFF; mem['h25CD]=8'hFF; mem['h25CE]=8'hFF; mem['h25CF]=8'hFF;
    mem['h25D0]=8'hFF; mem['h25D1]=8'hFF; mem['h25D2]=8'hFF; mem['h25D3]=8'hFF;
    mem['h25D4]=8'hFF; mem['h25D5]=8'hFF; mem['h25D6]=8'hFF; mem['h25D7]=8'hFF;
    mem['h25D8]=8'hFF; mem['h25D9]=8'hFF; mem['h25DA]=8'hFF; mem['h25DB]=8'hFF;
    mem['h25DC]=8'hFF; mem['h25DD]=8'hFF; mem['h25DE]=8'hFF; mem['h25DF]=8'hFF;
    mem['h25E0]=8'hFF; mem['h25E1]=8'hFF; mem['h25E2]=8'hFF; mem['h25E3]=8'hFF;
    mem['h25E4]=8'hFF; mem['h25E5]=8'hFF; mem['h25E6]=8'hFF; mem['h25E7]=8'hFF;
    mem['h25E8]=8'hFF; mem['h25E9]=8'hFF; mem['h25EA]=8'hFF; mem['h25EB]=8'hFF;
    mem['h25EC]=8'hFF; mem['h25ED]=8'hFF; mem['h25EE]=8'hFF; mem['h25EF]=8'hFF;
    mem['h25F0]=8'hFF; mem['h25F1]=8'hFF; mem['h25F2]=8'hFF; mem['h25F3]=8'hFF;
    mem['h25F4]=8'hFF; mem['h25F5]=8'hFF; mem['h25F6]=8'hFF; mem['h25F7]=8'hFF;
    mem['h25F8]=8'hFF; mem['h25F9]=8'hFF; mem['h25FA]=8'hFF; mem['h25FB]=8'hFF;
    mem['h25FC]=8'hFF; mem['h25FD]=8'hFF; mem['h25FE]=8'hFF; mem['h25FF]=8'hFF;
    mem['h2600]=8'hFF; mem['h2601]=8'hFF; mem['h2602]=8'hFF; mem['h2603]=8'hFF;
    mem['h2604]=8'hFF; mem['h2605]=8'hFF; mem['h2606]=8'hFF; mem['h2607]=8'hFF;
    mem['h2608]=8'hFF; mem['h2609]=8'hFF; mem['h260A]=8'hFF; mem['h260B]=8'hFF;
    mem['h260C]=8'hFF; mem['h260D]=8'hFF; mem['h260E]=8'hFF; mem['h260F]=8'hFF;
    mem['h2610]=8'hFF; mem['h2611]=8'hFF; mem['h2612]=8'hFF; mem['h2613]=8'hFF;
    mem['h2614]=8'hFF; mem['h2615]=8'hFF; mem['h2616]=8'hFF; mem['h2617]=8'hFF;
    mem['h2618]=8'hFF; mem['h2619]=8'hFF; mem['h261A]=8'hFF; mem['h261B]=8'hFF;
    mem['h261C]=8'hFF; mem['h261D]=8'hFF; mem['h261E]=8'hFF; mem['h261F]=8'hFF;
    mem['h2620]=8'hFF; mem['h2621]=8'hFF; mem['h2622]=8'hFF; mem['h2623]=8'hFF;
    mem['h2624]=8'hFF; mem['h2625]=8'hFF; mem['h2626]=8'hFF; mem['h2627]=8'hFF;
    mem['h2628]=8'hFF; mem['h2629]=8'hFF; mem['h262A]=8'hFF; mem['h262B]=8'hFF;
    mem['h262C]=8'hFF; mem['h262D]=8'hFF; mem['h262E]=8'hFF; mem['h262F]=8'hFF;
    mem['h2630]=8'hFF; mem['h2631]=8'hFF; mem['h2632]=8'hFF; mem['h2633]=8'hFF;
    mem['h2634]=8'hFF; mem['h2635]=8'hFF; mem['h2636]=8'hFF; mem['h2637]=8'hFF;
    mem['h2638]=8'hFF; mem['h2639]=8'hFF; mem['h263A]=8'hFF; mem['h263B]=8'hFF;
    mem['h263C]=8'hFF; mem['h263D]=8'hFF; mem['h263E]=8'hFF; mem['h263F]=8'hFF;
    mem['h2640]=8'hFF; mem['h2641]=8'hFF; mem['h2642]=8'hFF; mem['h2643]=8'hFF;
    mem['h2644]=8'hFF; mem['h2645]=8'hFF; mem['h2646]=8'hFF; mem['h2647]=8'hFF;
    mem['h2648]=8'hFF; mem['h2649]=8'hFF; mem['h264A]=8'hFF; mem['h264B]=8'hFF;
    mem['h264C]=8'hFF; mem['h264D]=8'hFF; mem['h264E]=8'hFF; mem['h264F]=8'hFF;
    mem['h2650]=8'hFF; mem['h2651]=8'hFF; mem['h2652]=8'hFF; mem['h2653]=8'hFF;
    mem['h2654]=8'hFF; mem['h2655]=8'hFF; mem['h2656]=8'hFF; mem['h2657]=8'hFF;
    mem['h2658]=8'hFF; mem['h2659]=8'hFF; mem['h265A]=8'hFF; mem['h265B]=8'hFF;
    mem['h265C]=8'hFF; mem['h265D]=8'hFF; mem['h265E]=8'hFF; mem['h265F]=8'hFF;
    mem['h2660]=8'hFF; mem['h2661]=8'hFF; mem['h2662]=8'hFF; mem['h2663]=8'hFF;
    mem['h2664]=8'hFF; mem['h2665]=8'hFF; mem['h2666]=8'hFF; mem['h2667]=8'hFF;
    mem['h2668]=8'hFF; mem['h2669]=8'hFF; mem['h266A]=8'hFF; mem['h266B]=8'hFF;
    mem['h266C]=8'hFF; mem['h266D]=8'hFF; mem['h266E]=8'hFF; mem['h266F]=8'hFF;
    mem['h2670]=8'hFF; mem['h2671]=8'hFF; mem['h2672]=8'hFF; mem['h2673]=8'hFF;
    mem['h2674]=8'hFF; mem['h2675]=8'hFF; mem['h2676]=8'hFF; mem['h2677]=8'hFF;
    mem['h2678]=8'hFF; mem['h2679]=8'hFF; mem['h267A]=8'hFF; mem['h267B]=8'hFF;
    mem['h267C]=8'hFF; mem['h267D]=8'hFF; mem['h267E]=8'hFF; mem['h267F]=8'hFF;
    mem['h2680]=8'hFF; mem['h2681]=8'hFF; mem['h2682]=8'hFF; mem['h2683]=8'hFF;
    mem['h2684]=8'hFF; mem['h2685]=8'hFF; mem['h2686]=8'hFF; mem['h2687]=8'hFF;
    mem['h2688]=8'hFF; mem['h2689]=8'hFF; mem['h268A]=8'hFF; mem['h268B]=8'hFF;
    mem['h268C]=8'hFF; mem['h268D]=8'hFF; mem['h268E]=8'hFF; mem['h268F]=8'hFF;
    mem['h2690]=8'hFF; mem['h2691]=8'hFF; mem['h2692]=8'hFF; mem['h2693]=8'hFF;
    mem['h2694]=8'hFF; mem['h2695]=8'hFF; mem['h2696]=8'hFF; mem['h2697]=8'hFF;
    mem['h2698]=8'hFF; mem['h2699]=8'hFF; mem['h269A]=8'hFF; mem['h269B]=8'hFF;
    mem['h269C]=8'hFF; mem['h269D]=8'hFF; mem['h269E]=8'hFF; mem['h269F]=8'hFF;
    mem['h26A0]=8'hFF; mem['h26A1]=8'hFF; mem['h26A2]=8'hFF; mem['h26A3]=8'hFF;
    mem['h26A4]=8'hFF; mem['h26A5]=8'hFF; mem['h26A6]=8'hFF; mem['h26A7]=8'hFF;
    mem['h26A8]=8'hFF; mem['h26A9]=8'hFF; mem['h26AA]=8'hFF; mem['h26AB]=8'hFF;
    mem['h26AC]=8'hFF; mem['h26AD]=8'hFF; mem['h26AE]=8'hFF; mem['h26AF]=8'hFF;
    mem['h26B0]=8'hFF; mem['h26B1]=8'hFF; mem['h26B2]=8'hFF; mem['h26B3]=8'hFF;
    mem['h26B4]=8'hFF; mem['h26B5]=8'hFF; mem['h26B6]=8'hFF; mem['h26B7]=8'hFF;
    mem['h26B8]=8'hFF; mem['h26B9]=8'hFF; mem['h26BA]=8'hFF; mem['h26BB]=8'hFF;
    mem['h26BC]=8'hFF; mem['h26BD]=8'hFF; mem['h26BE]=8'hFF; mem['h26BF]=8'hFF;
    mem['h26C0]=8'hFF; mem['h26C1]=8'hFF; mem['h26C2]=8'hFF; mem['h26C3]=8'hFF;
    mem['h26C4]=8'hFF; mem['h26C5]=8'hFF; mem['h26C6]=8'hFF; mem['h26C7]=8'hFF;
    mem['h26C8]=8'hFF; mem['h26C9]=8'hFF; mem['h26CA]=8'hFF; mem['h26CB]=8'hFF;
    mem['h26CC]=8'hFF; mem['h26CD]=8'hFF; mem['h26CE]=8'hFF; mem['h26CF]=8'hFF;
    mem['h26D0]=8'hFF; mem['h26D1]=8'hFF; mem['h26D2]=8'hFF; mem['h26D3]=8'hFF;
    mem['h26D4]=8'hFF; mem['h26D5]=8'hFF; mem['h26D6]=8'hFF; mem['h26D7]=8'hFF;
    mem['h26D8]=8'hFF; mem['h26D9]=8'hFF; mem['h26DA]=8'hFF; mem['h26DB]=8'hFF;
    mem['h26DC]=8'hFF; mem['h26DD]=8'hFF; mem['h26DE]=8'hFF; mem['h26DF]=8'hFF;
    mem['h26E0]=8'hFF; mem['h26E1]=8'hFF; mem['h26E2]=8'hFF; mem['h26E3]=8'hFF;
    mem['h26E4]=8'hFF; mem['h26E5]=8'hFF; mem['h26E6]=8'hFF; mem['h26E7]=8'hFF;
    mem['h26E8]=8'hFF; mem['h26E9]=8'hFF; mem['h26EA]=8'hFF; mem['h26EB]=8'hFF;
    mem['h26EC]=8'hFF; mem['h26ED]=8'hFF; mem['h26EE]=8'hFF; mem['h26EF]=8'hFF;
    mem['h26F0]=8'hFF; mem['h26F1]=8'hFF; mem['h26F2]=8'hFF; mem['h26F3]=8'hFF;
    mem['h26F4]=8'hFF; mem['h26F5]=8'hFF; mem['h26F6]=8'hFF; mem['h26F7]=8'hFF;
    mem['h26F8]=8'hFF; mem['h26F9]=8'hFF; mem['h26FA]=8'hFF; mem['h26FB]=8'hFF;
    mem['h26FC]=8'hFF; mem['h26FD]=8'hFF; mem['h26FE]=8'hFF; mem['h26FF]=8'hFF;
    mem['h2700]=8'hFF; mem['h2701]=8'hFF; mem['h2702]=8'hFF; mem['h2703]=8'hFF;
    mem['h2704]=8'hFF; mem['h2705]=8'hFF; mem['h2706]=8'hFF; mem['h2707]=8'hFF;
    mem['h2708]=8'hFF; mem['h2709]=8'hFF; mem['h270A]=8'hFF; mem['h270B]=8'hFF;
    mem['h270C]=8'hFF; mem['h270D]=8'hFF; mem['h270E]=8'hFF; mem['h270F]=8'hFF;
    mem['h2710]=8'hFF; mem['h2711]=8'hFF; mem['h2712]=8'hFF; mem['h2713]=8'hFF;
    mem['h2714]=8'hFF; mem['h2715]=8'hFF; mem['h2716]=8'hFF; mem['h2717]=8'hFF;
    mem['h2718]=8'hFF; mem['h2719]=8'hFF; mem['h271A]=8'hFF; mem['h271B]=8'hFF;
    mem['h271C]=8'hFF; mem['h271D]=8'hFF; mem['h271E]=8'hFF; mem['h271F]=8'hFF;
    mem['h2720]=8'hFF; mem['h2721]=8'hFF; mem['h2722]=8'hFF; mem['h2723]=8'hFF;
    mem['h2724]=8'hFF; mem['h2725]=8'hFF; mem['h2726]=8'hFF; mem['h2727]=8'hFF;
    mem['h2728]=8'hFF; mem['h2729]=8'hFF; mem['h272A]=8'hFF; mem['h272B]=8'hFF;
    mem['h272C]=8'hFF; mem['h272D]=8'hFF; mem['h272E]=8'hFF; mem['h272F]=8'hFF;
    mem['h2730]=8'hFF; mem['h2731]=8'hFF; mem['h2732]=8'hFF; mem['h2733]=8'hFF;
    mem['h2734]=8'hFF; mem['h2735]=8'hFF; mem['h2736]=8'hFF; mem['h2737]=8'hFF;
    mem['h2738]=8'hFF; mem['h2739]=8'hFF; mem['h273A]=8'hFF; mem['h273B]=8'hFF;
    mem['h273C]=8'hFF; mem['h273D]=8'hFF; mem['h273E]=8'hFF; mem['h273F]=8'hFF;
    mem['h2740]=8'hFF; mem['h2741]=8'hFF; mem['h2742]=8'hFF; mem['h2743]=8'hFF;
    mem['h2744]=8'hFF; mem['h2745]=8'hFF; mem['h2746]=8'hFF; mem['h2747]=8'hFF;
    mem['h2748]=8'hFF; mem['h2749]=8'hFF; mem['h274A]=8'hFF; mem['h274B]=8'hFF;
    mem['h274C]=8'hFF; mem['h274D]=8'hFF; mem['h274E]=8'hFF; mem['h274F]=8'hFF;
    mem['h2750]=8'hFF; mem['h2751]=8'hFF; mem['h2752]=8'hFF; mem['h2753]=8'hFF;
    mem['h2754]=8'hFF; mem['h2755]=8'hFF; mem['h2756]=8'hFF; mem['h2757]=8'hFF;
    mem['h2758]=8'hFF; mem['h2759]=8'hFF; mem['h275A]=8'hFF; mem['h275B]=8'hFF;
    mem['h275C]=8'hFF; mem['h275D]=8'hFF; mem['h275E]=8'hFF; mem['h275F]=8'hFF;
    mem['h2760]=8'hFF; mem['h2761]=8'hFF; mem['h2762]=8'hFF; mem['h2763]=8'hFF;
    mem['h2764]=8'hFF; mem['h2765]=8'hFF; mem['h2766]=8'hFF; mem['h2767]=8'hFF;
    mem['h2768]=8'hFF; mem['h2769]=8'hFF; mem['h276A]=8'hFF; mem['h276B]=8'hFF;
    mem['h276C]=8'hFF; mem['h276D]=8'hFF; mem['h276E]=8'hFF; mem['h276F]=8'hFF;
    mem['h2770]=8'hFF; mem['h2771]=8'hFF; mem['h2772]=8'hFF; mem['h2773]=8'hFF;
    mem['h2774]=8'hFF; mem['h2775]=8'hFF; mem['h2776]=8'hFF; mem['h2777]=8'hFF;
    mem['h2778]=8'hFF; mem['h2779]=8'hFF; mem['h277A]=8'hFF; mem['h277B]=8'hFF;
    mem['h277C]=8'hFF; mem['h277D]=8'hFF; mem['h277E]=8'hFF; mem['h277F]=8'hFF;
    mem['h2780]=8'hFF; mem['h2781]=8'hFF; mem['h2782]=8'hFF; mem['h2783]=8'hFF;
    mem['h2784]=8'hFF; mem['h2785]=8'hFF; mem['h2786]=8'hFF; mem['h2787]=8'hFF;
    mem['h2788]=8'hFF; mem['h2789]=8'hFF; mem['h278A]=8'hFF; mem['h278B]=8'hFF;
    mem['h278C]=8'hFF; mem['h278D]=8'hFF; mem['h278E]=8'hFF; mem['h278F]=8'hFF;
    mem['h2790]=8'hFF; mem['h2791]=8'hFF; mem['h2792]=8'hFF; mem['h2793]=8'hFF;
    mem['h2794]=8'hFF; mem['h2795]=8'hFF; mem['h2796]=8'hFF; mem['h2797]=8'hFF;
    mem['h2798]=8'hFF; mem['h2799]=8'hFF; mem['h279A]=8'hFF; mem['h279B]=8'hFF;
    mem['h279C]=8'hFF; mem['h279D]=8'hFF; mem['h279E]=8'hFF; mem['h279F]=8'hFF;
    mem['h27A0]=8'hFF; mem['h27A1]=8'hFF; mem['h27A2]=8'hFF; mem['h27A3]=8'hFF;
    mem['h27A4]=8'hFF; mem['h27A5]=8'hFF; mem['h27A6]=8'hFF; mem['h27A7]=8'hFF;
    mem['h27A8]=8'hFF; mem['h27A9]=8'hFF; mem['h27AA]=8'hFF; mem['h27AB]=8'hFF;
    mem['h27AC]=8'hFF; mem['h27AD]=8'hFF; mem['h27AE]=8'hFF; mem['h27AF]=8'hFF;
    mem['h27B0]=8'hFF; mem['h27B1]=8'hFF; mem['h27B2]=8'hFF; mem['h27B3]=8'hFF;
    mem['h27B4]=8'hFF; mem['h27B5]=8'hFF; mem['h27B6]=8'hFF; mem['h27B7]=8'hFF;
    mem['h27B8]=8'hFF; mem['h27B9]=8'hFF; mem['h27BA]=8'hFF; mem['h27BB]=8'hFF;
    mem['h27BC]=8'hFF; mem['h27BD]=8'hFF; mem['h27BE]=8'hFF; mem['h27BF]=8'hFF;
    mem['h27C0]=8'hFF; mem['h27C1]=8'hFF; mem['h27C2]=8'hFF; mem['h27C3]=8'hFF;
    mem['h27C4]=8'hFF; mem['h27C5]=8'hFF; mem['h27C6]=8'hFF; mem['h27C7]=8'hFF;
    mem['h27C8]=8'hFF; mem['h27C9]=8'hFF; mem['h27CA]=8'hFF; mem['h27CB]=8'hFF;
    mem['h27CC]=8'hFF; mem['h27CD]=8'hFF; mem['h27CE]=8'hFF; mem['h27CF]=8'hFF;
    mem['h27D0]=8'hFF; mem['h27D1]=8'hFF; mem['h27D2]=8'hFF; mem['h27D3]=8'hFF;
    mem['h27D4]=8'hFF; mem['h27D5]=8'hFF; mem['h27D6]=8'hFF; mem['h27D7]=8'hFF;
    mem['h27D8]=8'hFF; mem['h27D9]=8'hFF; mem['h27DA]=8'hFF; mem['h27DB]=8'hFF;
    mem['h27DC]=8'hFF; mem['h27DD]=8'hFF; mem['h27DE]=8'hFF; mem['h27DF]=8'hFF;
    mem['h27E0]=8'hFF; mem['h27E1]=8'hFF; mem['h27E2]=8'hFF; mem['h27E3]=8'hFF;
    mem['h27E4]=8'hFF; mem['h27E5]=8'hFF; mem['h27E6]=8'hFF; mem['h27E7]=8'hFF;
    mem['h27E8]=8'hFF; mem['h27E9]=8'hFF; mem['h27EA]=8'hFF; mem['h27EB]=8'hFF;
    mem['h27EC]=8'hFF; mem['h27ED]=8'hFF; mem['h27EE]=8'hFF; mem['h27EF]=8'hFF;
    mem['h27F0]=8'hFF; mem['h27F1]=8'hFF; mem['h27F2]=8'hFF; mem['h27F3]=8'hFF;
    mem['h27F4]=8'hFF; mem['h27F5]=8'hFF; mem['h27F6]=8'hFF; mem['h27F7]=8'hFF;
    mem['h27F8]=8'hFF; mem['h27F9]=8'hFF; mem['h27FA]=8'hFF; mem['h27FB]=8'hFF;
    mem['h27FC]=8'hFF; mem['h27FD]=8'hFF; mem['h27FE]=8'hFF; mem['h27FF]=8'hFF;
    mem['h2800]=8'hFF; mem['h2801]=8'hFF; mem['h2802]=8'hFF; mem['h2803]=8'hFF;
    mem['h2804]=8'hFF; mem['h2805]=8'hFF; mem['h2806]=8'hFF; mem['h2807]=8'hFF;
    mem['h2808]=8'hFF; mem['h2809]=8'hFF; mem['h280A]=8'hFF; mem['h280B]=8'hFF;
    mem['h280C]=8'hFF; mem['h280D]=8'hFF; mem['h280E]=8'hFF; mem['h280F]=8'hFF;
    mem['h2810]=8'hFF; mem['h2811]=8'hFF; mem['h2812]=8'hFF; mem['h2813]=8'hFF;
    mem['h2814]=8'hFF; mem['h2815]=8'hFF; mem['h2816]=8'hFF; mem['h2817]=8'hFF;
    mem['h2818]=8'hFF; mem['h2819]=8'hFF; mem['h281A]=8'hFF; mem['h281B]=8'hFF;
    mem['h281C]=8'hFF; mem['h281D]=8'hFF; mem['h281E]=8'hFF; mem['h281F]=8'hFF;
    mem['h2820]=8'hFF; mem['h2821]=8'hFF; mem['h2822]=8'hFF; mem['h2823]=8'hFF;
    mem['h2824]=8'hFF; mem['h2825]=8'hFF; mem['h2826]=8'hFF; mem['h2827]=8'hFF;
    mem['h2828]=8'hFF; mem['h2829]=8'hFF; mem['h282A]=8'hFF; mem['h282B]=8'hFF;
    mem['h282C]=8'hFF; mem['h282D]=8'hFF; mem['h282E]=8'hFF; mem['h282F]=8'hFF;
    mem['h2830]=8'hFF; mem['h2831]=8'hFF; mem['h2832]=8'hFF; mem['h2833]=8'hFF;
    mem['h2834]=8'hFF; mem['h2835]=8'hFF; mem['h2836]=8'hFF; mem['h2837]=8'hFF;
    mem['h2838]=8'hFF; mem['h2839]=8'hFF; mem['h283A]=8'hFF; mem['h283B]=8'hFF;
    mem['h283C]=8'hFF; mem['h283D]=8'hFF; mem['h283E]=8'hFF; mem['h283F]=8'hFF;
    mem['h2840]=8'hFF; mem['h2841]=8'hFF; mem['h2842]=8'hFF; mem['h2843]=8'hFF;
    mem['h2844]=8'hFF; mem['h2845]=8'hFF; mem['h2846]=8'hFF; mem['h2847]=8'hFF;
    mem['h2848]=8'hFF; mem['h2849]=8'hFF; mem['h284A]=8'hFF; mem['h284B]=8'hFF;
    mem['h284C]=8'hFF; mem['h284D]=8'hFF; mem['h284E]=8'hFF; mem['h284F]=8'hFF;
    mem['h2850]=8'hFF; mem['h2851]=8'hFF; mem['h2852]=8'hFF; mem['h2853]=8'hFF;
    mem['h2854]=8'hFF; mem['h2855]=8'hFF; mem['h2856]=8'hFF; mem['h2857]=8'hFF;
    mem['h2858]=8'hFF; mem['h2859]=8'hFF; mem['h285A]=8'hFF; mem['h285B]=8'hFF;
    mem['h285C]=8'hFF; mem['h285D]=8'hFF; mem['h285E]=8'hFF; mem['h285F]=8'hFF;
    mem['h2860]=8'hFF; mem['h2861]=8'hFF; mem['h2862]=8'hFF; mem['h2863]=8'hFF;
    mem['h2864]=8'hFF; mem['h2865]=8'hFF; mem['h2866]=8'hFF; mem['h2867]=8'hFF;
    mem['h2868]=8'hFF; mem['h2869]=8'hFF; mem['h286A]=8'hFF; mem['h286B]=8'hFF;
    mem['h286C]=8'hFF; mem['h286D]=8'hFF; mem['h286E]=8'hFF; mem['h286F]=8'hFF;
    mem['h2870]=8'hFF; mem['h2871]=8'hFF; mem['h2872]=8'hFF; mem['h2873]=8'hFF;
    mem['h2874]=8'hFF; mem['h2875]=8'hFF; mem['h2876]=8'hFF; mem['h2877]=8'hFF;
    mem['h2878]=8'hFF; mem['h2879]=8'hFF; mem['h287A]=8'hFF; mem['h287B]=8'hFF;
    mem['h287C]=8'hFF; mem['h287D]=8'hFF; mem['h287E]=8'hFF; mem['h287F]=8'hFF;
    mem['h2880]=8'hFF; mem['h2881]=8'hFF; mem['h2882]=8'hFF; mem['h2883]=8'hFF;
    mem['h2884]=8'hFF; mem['h2885]=8'hFF; mem['h2886]=8'hFF; mem['h2887]=8'hFF;
    mem['h2888]=8'hFF; mem['h2889]=8'hFF; mem['h288A]=8'hFF; mem['h288B]=8'hFF;
    mem['h288C]=8'hFF; mem['h288D]=8'hFF; mem['h288E]=8'hFF; mem['h288F]=8'hFF;
    mem['h2890]=8'hFF; mem['h2891]=8'hFF; mem['h2892]=8'hFF; mem['h2893]=8'hFF;
    mem['h2894]=8'hFF; mem['h2895]=8'hFF; mem['h2896]=8'hFF; mem['h2897]=8'hFF;
    mem['h2898]=8'hFF; mem['h2899]=8'hFF; mem['h289A]=8'hFF; mem['h289B]=8'hFF;
    mem['h289C]=8'hFF; mem['h289D]=8'hFF; mem['h289E]=8'hFF; mem['h289F]=8'hFF;
    mem['h28A0]=8'hFF; mem['h28A1]=8'hFF; mem['h28A2]=8'hFF; mem['h28A3]=8'hFF;
    mem['h28A4]=8'hFF; mem['h28A5]=8'hFF; mem['h28A6]=8'hFF; mem['h28A7]=8'hFF;
    mem['h28A8]=8'hFF; mem['h28A9]=8'hFF; mem['h28AA]=8'hFF; mem['h28AB]=8'hFF;
    mem['h28AC]=8'hFF; mem['h28AD]=8'hFF; mem['h28AE]=8'hFF; mem['h28AF]=8'hFF;
    mem['h28B0]=8'hFF; mem['h28B1]=8'hFF; mem['h28B2]=8'hFF; mem['h28B3]=8'hFF;
    mem['h28B4]=8'hFF; mem['h28B5]=8'hFF; mem['h28B6]=8'hFF; mem['h28B7]=8'hFF;
    mem['h28B8]=8'hFF; mem['h28B9]=8'hFF; mem['h28BA]=8'hFF; mem['h28BB]=8'hFF;
    mem['h28BC]=8'hFF; mem['h28BD]=8'hFF; mem['h28BE]=8'hFF; mem['h28BF]=8'hFF;
    mem['h28C0]=8'hFF; mem['h28C1]=8'hFF; mem['h28C2]=8'hFF; mem['h28C3]=8'hFF;
    mem['h28C4]=8'hFF; mem['h28C5]=8'hFF; mem['h28C6]=8'hFF; mem['h28C7]=8'hFF;
    mem['h28C8]=8'hFF; mem['h28C9]=8'hFF; mem['h28CA]=8'hFF; mem['h28CB]=8'hFF;
    mem['h28CC]=8'hFF; mem['h28CD]=8'hFF; mem['h28CE]=8'hFF; mem['h28CF]=8'hFF;
    mem['h28D0]=8'hFF; mem['h28D1]=8'hFF; mem['h28D2]=8'hFF; mem['h28D3]=8'hFF;
    mem['h28D4]=8'hFF; mem['h28D5]=8'hFF; mem['h28D6]=8'hFF; mem['h28D7]=8'hFF;
    mem['h28D8]=8'hFF; mem['h28D9]=8'hFF; mem['h28DA]=8'hFF; mem['h28DB]=8'hFF;
    mem['h28DC]=8'hFF; mem['h28DD]=8'hFF; mem['h28DE]=8'hFF; mem['h28DF]=8'hFF;
    mem['h28E0]=8'hFF; mem['h28E1]=8'hFF; mem['h28E2]=8'hFF; mem['h28E3]=8'hFF;
    mem['h28E4]=8'hFF; mem['h28E5]=8'hFF; mem['h28E6]=8'hFF; mem['h28E7]=8'hFF;
    mem['h28E8]=8'hFF; mem['h28E9]=8'hFF; mem['h28EA]=8'hFF; mem['h28EB]=8'hFF;
    mem['h28EC]=8'hFF; mem['h28ED]=8'hFF; mem['h28EE]=8'hFF; mem['h28EF]=8'hFF;
    mem['h28F0]=8'hFF; mem['h28F1]=8'hFF; mem['h28F2]=8'hFF; mem['h28F3]=8'hFF;
    mem['h28F4]=8'hFF; mem['h28F5]=8'hFF; mem['h28F6]=8'hFF; mem['h28F7]=8'hFF;
    mem['h28F8]=8'hFF; mem['h28F9]=8'hFF; mem['h28FA]=8'hFF; mem['h28FB]=8'hFF;
    mem['h28FC]=8'hFF; mem['h28FD]=8'hFF; mem['h28FE]=8'hFF; mem['h28FF]=8'hFF;
    mem['h2900]=8'hFF; mem['h2901]=8'hFF; mem['h2902]=8'hFF; mem['h2903]=8'hFF;
    mem['h2904]=8'hFF; mem['h2905]=8'hFF; mem['h2906]=8'hFF; mem['h2907]=8'hFF;
    mem['h2908]=8'hFF; mem['h2909]=8'hFF; mem['h290A]=8'hFF; mem['h290B]=8'hFF;
    mem['h290C]=8'hFF; mem['h290D]=8'hFF; mem['h290E]=8'hFF; mem['h290F]=8'hFF;
    mem['h2910]=8'hFF; mem['h2911]=8'hFF; mem['h2912]=8'hFF; mem['h2913]=8'hFF;
    mem['h2914]=8'hFF; mem['h2915]=8'hFF; mem['h2916]=8'hFF; mem['h2917]=8'hFF;
    mem['h2918]=8'hFF; mem['h2919]=8'hFF; mem['h291A]=8'hFF; mem['h291B]=8'hFF;
    mem['h291C]=8'hFF; mem['h291D]=8'hFF; mem['h291E]=8'hFF; mem['h291F]=8'hFF;
    mem['h2920]=8'hFF; mem['h2921]=8'hFF; mem['h2922]=8'hFF; mem['h2923]=8'hFF;
    mem['h2924]=8'hFF; mem['h2925]=8'hFF; mem['h2926]=8'hFF; mem['h2927]=8'hFF;
    mem['h2928]=8'hFF; mem['h2929]=8'hFF; mem['h292A]=8'hFF; mem['h292B]=8'hFF;
    mem['h292C]=8'hFF; mem['h292D]=8'hFF; mem['h292E]=8'hFF; mem['h292F]=8'hFF;
    mem['h2930]=8'hFF; mem['h2931]=8'hFF; mem['h2932]=8'hFF; mem['h2933]=8'hFF;
    mem['h2934]=8'hFF; mem['h2935]=8'hFF; mem['h2936]=8'hFF; mem['h2937]=8'hFF;
    mem['h2938]=8'hFF; mem['h2939]=8'hFF; mem['h293A]=8'hFF; mem['h293B]=8'hFF;
    mem['h293C]=8'hFF; mem['h293D]=8'hFF; mem['h293E]=8'hFF; mem['h293F]=8'hFF;
    mem['h2940]=8'hFF; mem['h2941]=8'hFF; mem['h2942]=8'hFF; mem['h2943]=8'hFF;
    mem['h2944]=8'hFF; mem['h2945]=8'hFF; mem['h2946]=8'hFF; mem['h2947]=8'hFF;
    mem['h2948]=8'hFF; mem['h2949]=8'hFF; mem['h294A]=8'hFF; mem['h294B]=8'hFF;
    mem['h294C]=8'hFF; mem['h294D]=8'hFF; mem['h294E]=8'hFF; mem['h294F]=8'hFF;
    mem['h2950]=8'hFF; mem['h2951]=8'hFF; mem['h2952]=8'hFF; mem['h2953]=8'hFF;
    mem['h2954]=8'hFF; mem['h2955]=8'hFF; mem['h2956]=8'hFF; mem['h2957]=8'hFF;
    mem['h2958]=8'hFF; mem['h2959]=8'hFF; mem['h295A]=8'hFF; mem['h295B]=8'hFF;
    mem['h295C]=8'hFF; mem['h295D]=8'hFF; mem['h295E]=8'hFF; mem['h295F]=8'hFF;
    mem['h2960]=8'hFF; mem['h2961]=8'hFF; mem['h2962]=8'hFF; mem['h2963]=8'hFF;
    mem['h2964]=8'hFF; mem['h2965]=8'hFF; mem['h2966]=8'hFF; mem['h2967]=8'hFF;
    mem['h2968]=8'hFF; mem['h2969]=8'hFF; mem['h296A]=8'hFF; mem['h296B]=8'hFF;
    mem['h296C]=8'hFF; mem['h296D]=8'hFF; mem['h296E]=8'hFF; mem['h296F]=8'hFF;
    mem['h2970]=8'hFF; mem['h2971]=8'hFF; mem['h2972]=8'hFF; mem['h2973]=8'hFF;
    mem['h2974]=8'hFF; mem['h2975]=8'hFF; mem['h2976]=8'hFF; mem['h2977]=8'hFF;
    mem['h2978]=8'hFF; mem['h2979]=8'hFF; mem['h297A]=8'hFF; mem['h297B]=8'hFF;
    mem['h297C]=8'hFF; mem['h297D]=8'hFF; mem['h297E]=8'hFF; mem['h297F]=8'hFF;
    mem['h2980]=8'hFF; mem['h2981]=8'hFF; mem['h2982]=8'hFF; mem['h2983]=8'hFF;
    mem['h2984]=8'hFF; mem['h2985]=8'hFF; mem['h2986]=8'hFF; mem['h2987]=8'hFF;
    mem['h2988]=8'hFF; mem['h2989]=8'hFF; mem['h298A]=8'hFF; mem['h298B]=8'hFF;
    mem['h298C]=8'hFF; mem['h298D]=8'hFF; mem['h298E]=8'hFF; mem['h298F]=8'hFF;
    mem['h2990]=8'hFF; mem['h2991]=8'hFF; mem['h2992]=8'hFF; mem['h2993]=8'hFF;
    mem['h2994]=8'hFF; mem['h2995]=8'hFF; mem['h2996]=8'hFF; mem['h2997]=8'hFF;
    mem['h2998]=8'hFF; mem['h2999]=8'hFF; mem['h299A]=8'hFF; mem['h299B]=8'hFF;
    mem['h299C]=8'hFF; mem['h299D]=8'hFF; mem['h299E]=8'hFF; mem['h299F]=8'hFF;
    mem['h29A0]=8'hFF; mem['h29A1]=8'hFF; mem['h29A2]=8'hFF; mem['h29A3]=8'hFF;
    mem['h29A4]=8'hFF; mem['h29A5]=8'hFF; mem['h29A6]=8'hFF; mem['h29A7]=8'hFF;
    mem['h29A8]=8'hFF; mem['h29A9]=8'hFF; mem['h29AA]=8'hFF; mem['h29AB]=8'hFF;
    mem['h29AC]=8'hFF; mem['h29AD]=8'hFF; mem['h29AE]=8'hFF; mem['h29AF]=8'hFF;
    mem['h29B0]=8'hFF; mem['h29B1]=8'hFF; mem['h29B2]=8'hFF; mem['h29B3]=8'hFF;
    mem['h29B4]=8'hFF; mem['h29B5]=8'hFF; mem['h29B6]=8'hFF; mem['h29B7]=8'hFF;
    mem['h29B8]=8'hFF; mem['h29B9]=8'hFF; mem['h29BA]=8'hFF; mem['h29BB]=8'hFF;
    mem['h29BC]=8'hFF; mem['h29BD]=8'hFF; mem['h29BE]=8'hFF; mem['h29BF]=8'hFF;
    mem['h29C0]=8'hFF; mem['h29C1]=8'hFF; mem['h29C2]=8'hFF; mem['h29C3]=8'hFF;
    mem['h29C4]=8'hFF; mem['h29C5]=8'hFF; mem['h29C6]=8'hFF; mem['h29C7]=8'hFF;
    mem['h29C8]=8'hFF; mem['h29C9]=8'hFF; mem['h29CA]=8'hFF; mem['h29CB]=8'hFF;
    mem['h29CC]=8'hFF; mem['h29CD]=8'hFF; mem['h29CE]=8'hFF; mem['h29CF]=8'hFF;
    mem['h29D0]=8'hFF; mem['h29D1]=8'hFF; mem['h29D2]=8'hFF; mem['h29D3]=8'hFF;
    mem['h29D4]=8'hFF; mem['h29D5]=8'hFF; mem['h29D6]=8'hFF; mem['h29D7]=8'hFF;
    mem['h29D8]=8'hFF; mem['h29D9]=8'hFF; mem['h29DA]=8'hFF; mem['h29DB]=8'hFF;
    mem['h29DC]=8'hFF; mem['h29DD]=8'hFF; mem['h29DE]=8'hFF; mem['h29DF]=8'hFF;
    mem['h29E0]=8'hFF; mem['h29E1]=8'hFF; mem['h29E2]=8'hFF; mem['h29E3]=8'hFF;
    mem['h29E4]=8'hFF; mem['h29E5]=8'hFF; mem['h29E6]=8'hFF; mem['h29E7]=8'hFF;
    mem['h29E8]=8'hFF; mem['h29E9]=8'hFF; mem['h29EA]=8'hFF; mem['h29EB]=8'hFF;
    mem['h29EC]=8'hFF; mem['h29ED]=8'hFF; mem['h29EE]=8'hFF; mem['h29EF]=8'hFF;
    mem['h29F0]=8'hFF; mem['h29F1]=8'hFF; mem['h29F2]=8'hFF; mem['h29F3]=8'hFF;
    mem['h29F4]=8'hFF; mem['h29F5]=8'hFF; mem['h29F6]=8'hFF; mem['h29F7]=8'hFF;
    mem['h29F8]=8'hFF; mem['h29F9]=8'hFF; mem['h29FA]=8'hFF; mem['h29FB]=8'hFF;
    mem['h29FC]=8'hFF; mem['h29FD]=8'hFF; mem['h29FE]=8'hFF; mem['h29FF]=8'hFF;
    mem['h2A00]=8'hFF; mem['h2A01]=8'hFF; mem['h2A02]=8'hFF; mem['h2A03]=8'hFF;
    mem['h2A04]=8'hFF; mem['h2A05]=8'hFF; mem['h2A06]=8'hFF; mem['h2A07]=8'hFF;
    mem['h2A08]=8'hFF; mem['h2A09]=8'hFF; mem['h2A0A]=8'hFF; mem['h2A0B]=8'hFF;
    mem['h2A0C]=8'hFF; mem['h2A0D]=8'hFF; mem['h2A0E]=8'hFF; mem['h2A0F]=8'hFF;
    mem['h2A10]=8'hFF; mem['h2A11]=8'hFF; mem['h2A12]=8'hFF; mem['h2A13]=8'hFF;
    mem['h2A14]=8'hFF; mem['h2A15]=8'hFF; mem['h2A16]=8'hFF; mem['h2A17]=8'hFF;
    mem['h2A18]=8'hFF; mem['h2A19]=8'hFF; mem['h2A1A]=8'hFF; mem['h2A1B]=8'hFF;
    mem['h2A1C]=8'hFF; mem['h2A1D]=8'hFF; mem['h2A1E]=8'hFF; mem['h2A1F]=8'hFF;
    mem['h2A20]=8'hFF; mem['h2A21]=8'hFF; mem['h2A22]=8'hFF; mem['h2A23]=8'hFF;
    mem['h2A24]=8'hFF; mem['h2A25]=8'hFF; mem['h2A26]=8'hFF; mem['h2A27]=8'hFF;
    mem['h2A28]=8'hFF; mem['h2A29]=8'hFF; mem['h2A2A]=8'hFF; mem['h2A2B]=8'hFF;
    mem['h2A2C]=8'hFF; mem['h2A2D]=8'hFF; mem['h2A2E]=8'hFF; mem['h2A2F]=8'hFF;
    mem['h2A30]=8'hFF; mem['h2A31]=8'hFF; mem['h2A32]=8'hFF; mem['h2A33]=8'hFF;
    mem['h2A34]=8'hFF; mem['h2A35]=8'hFF; mem['h2A36]=8'hFF; mem['h2A37]=8'hFF;
    mem['h2A38]=8'hFF; mem['h2A39]=8'hFF; mem['h2A3A]=8'hFF; mem['h2A3B]=8'hFF;
    mem['h2A3C]=8'hFF; mem['h2A3D]=8'hFF; mem['h2A3E]=8'hFF; mem['h2A3F]=8'hFF;
    mem['h2A40]=8'hFF; mem['h2A41]=8'hFF; mem['h2A42]=8'hFF; mem['h2A43]=8'hFF;
    mem['h2A44]=8'hFF; mem['h2A45]=8'hFF; mem['h2A46]=8'hFF; mem['h2A47]=8'hFF;
    mem['h2A48]=8'hFF; mem['h2A49]=8'hFF; mem['h2A4A]=8'hFF; mem['h2A4B]=8'hFF;
    mem['h2A4C]=8'hFF; mem['h2A4D]=8'hFF; mem['h2A4E]=8'hFF; mem['h2A4F]=8'hFF;
    mem['h2A50]=8'hFF; mem['h2A51]=8'hFF; mem['h2A52]=8'hFF; mem['h2A53]=8'hFF;
    mem['h2A54]=8'hFF; mem['h2A55]=8'hFF; mem['h2A56]=8'hFF; mem['h2A57]=8'hFF;
    mem['h2A58]=8'hFF; mem['h2A59]=8'hFF; mem['h2A5A]=8'hFF; mem['h2A5B]=8'hFF;
    mem['h2A5C]=8'hFF; mem['h2A5D]=8'hFF; mem['h2A5E]=8'hFF; mem['h2A5F]=8'hFF;
    mem['h2A60]=8'hFF; mem['h2A61]=8'hFF; mem['h2A62]=8'hFF; mem['h2A63]=8'hFF;
    mem['h2A64]=8'hFF; mem['h2A65]=8'hFF; mem['h2A66]=8'hFF; mem['h2A67]=8'hFF;
    mem['h2A68]=8'hFF; mem['h2A69]=8'hFF; mem['h2A6A]=8'hFF; mem['h2A6B]=8'hFF;
    mem['h2A6C]=8'hFF; mem['h2A6D]=8'hFF; mem['h2A6E]=8'hFF; mem['h2A6F]=8'hFF;
    mem['h2A70]=8'hFF; mem['h2A71]=8'hFF; mem['h2A72]=8'hFF; mem['h2A73]=8'hFF;
    mem['h2A74]=8'hFF; mem['h2A75]=8'hFF; mem['h2A76]=8'hFF; mem['h2A77]=8'hFF;
    mem['h2A78]=8'hFF; mem['h2A79]=8'hFF; mem['h2A7A]=8'hFF; mem['h2A7B]=8'hFF;
    mem['h2A7C]=8'hFF; mem['h2A7D]=8'hFF; mem['h2A7E]=8'hFF; mem['h2A7F]=8'hFF;
    mem['h2A80]=8'hFF; mem['h2A81]=8'hFF; mem['h2A82]=8'hFF; mem['h2A83]=8'hFF;
    mem['h2A84]=8'hFF; mem['h2A85]=8'hFF; mem['h2A86]=8'hFF; mem['h2A87]=8'hFF;
    mem['h2A88]=8'hFF; mem['h2A89]=8'hFF; mem['h2A8A]=8'hFF; mem['h2A8B]=8'hFF;
    mem['h2A8C]=8'hFF; mem['h2A8D]=8'hFF; mem['h2A8E]=8'hFF; mem['h2A8F]=8'hFF;
    mem['h2A90]=8'hFF; mem['h2A91]=8'hFF; mem['h2A92]=8'hFF; mem['h2A93]=8'hFF;
    mem['h2A94]=8'hFF; mem['h2A95]=8'hFF; mem['h2A96]=8'hFF; mem['h2A97]=8'hFF;
    mem['h2A98]=8'hFF; mem['h2A99]=8'hFF; mem['h2A9A]=8'hFF; mem['h2A9B]=8'hFF;
    mem['h2A9C]=8'hFF; mem['h2A9D]=8'hFF; mem['h2A9E]=8'hFF; mem['h2A9F]=8'hFF;
    mem['h2AA0]=8'hFF; mem['h2AA1]=8'hFF; mem['h2AA2]=8'hFF; mem['h2AA3]=8'hFF;
    mem['h2AA4]=8'hFF; mem['h2AA5]=8'hFF; mem['h2AA6]=8'hFF; mem['h2AA7]=8'hFF;
    mem['h2AA8]=8'hFF; mem['h2AA9]=8'hFF; mem['h2AAA]=8'hFF; mem['h2AAB]=8'hFF;
    mem['h2AAC]=8'hFF; mem['h2AAD]=8'hFF; mem['h2AAE]=8'hFF; mem['h2AAF]=8'hFF;
    mem['h2AB0]=8'hFF; mem['h2AB1]=8'hFF; mem['h2AB2]=8'hFF; mem['h2AB3]=8'hFF;
    mem['h2AB4]=8'hFF; mem['h2AB5]=8'hFF; mem['h2AB6]=8'hFF; mem['h2AB7]=8'hFF;
    mem['h2AB8]=8'hFF; mem['h2AB9]=8'hFF; mem['h2ABA]=8'hFF; mem['h2ABB]=8'hFF;
    mem['h2ABC]=8'hFF; mem['h2ABD]=8'hFF; mem['h2ABE]=8'hFF; mem['h2ABF]=8'hFF;
    mem['h2AC0]=8'hFF; mem['h2AC1]=8'hFF; mem['h2AC2]=8'hFF; mem['h2AC3]=8'hFF;
    mem['h2AC4]=8'hFF; mem['h2AC5]=8'hFF; mem['h2AC6]=8'hFF; mem['h2AC7]=8'hFF;
    mem['h2AC8]=8'hFF; mem['h2AC9]=8'hFF; mem['h2ACA]=8'hFF; mem['h2ACB]=8'hFF;
    mem['h2ACC]=8'hFF; mem['h2ACD]=8'hFF; mem['h2ACE]=8'hFF; mem['h2ACF]=8'hFF;
    mem['h2AD0]=8'hFF; mem['h2AD1]=8'hFF; mem['h2AD2]=8'hFF; mem['h2AD3]=8'hFF;
    mem['h2AD4]=8'hFF; mem['h2AD5]=8'hFF; mem['h2AD6]=8'hFF; mem['h2AD7]=8'hFF;
    mem['h2AD8]=8'hFF; mem['h2AD9]=8'hFF; mem['h2ADA]=8'hFF; mem['h2ADB]=8'hFF;
    mem['h2ADC]=8'hFF; mem['h2ADD]=8'hFF; mem['h2ADE]=8'hFF; mem['h2ADF]=8'hFF;
    mem['h2AE0]=8'hFF; mem['h2AE1]=8'hFF; mem['h2AE2]=8'hFF; mem['h2AE3]=8'hFF;
    mem['h2AE4]=8'hFF; mem['h2AE5]=8'hFF; mem['h2AE6]=8'hFF; mem['h2AE7]=8'hFF;
    mem['h2AE8]=8'hFF; mem['h2AE9]=8'hFF; mem['h2AEA]=8'hFF; mem['h2AEB]=8'hFF;
    mem['h2AEC]=8'hFF; mem['h2AED]=8'hFF; mem['h2AEE]=8'hFF; mem['h2AEF]=8'hFF;
    mem['h2AF0]=8'hFF; mem['h2AF1]=8'hFF; mem['h2AF2]=8'hFF; mem['h2AF3]=8'hFF;
    mem['h2AF4]=8'hFF; mem['h2AF5]=8'hFF; mem['h2AF6]=8'hFF; mem['h2AF7]=8'hFF;
    mem['h2AF8]=8'hFF; mem['h2AF9]=8'hFF; mem['h2AFA]=8'hFF; mem['h2AFB]=8'hFF;
    mem['h2AFC]=8'hFF; mem['h2AFD]=8'hFF; mem['h2AFE]=8'hFF; mem['h2AFF]=8'hFF;
    mem['h2B00]=8'hFF; mem['h2B01]=8'hFF; mem['h2B02]=8'hFF; mem['h2B03]=8'hFF;
    mem['h2B04]=8'hFF; mem['h2B05]=8'hFF; mem['h2B06]=8'hFF; mem['h2B07]=8'hFF;
    mem['h2B08]=8'hFF; mem['h2B09]=8'hFF; mem['h2B0A]=8'hFF; mem['h2B0B]=8'hFF;
    mem['h2B0C]=8'hFF; mem['h2B0D]=8'hFF; mem['h2B0E]=8'hFF; mem['h2B0F]=8'hFF;
    mem['h2B10]=8'hFF; mem['h2B11]=8'hFF; mem['h2B12]=8'hFF; mem['h2B13]=8'hFF;
    mem['h2B14]=8'hFF; mem['h2B15]=8'hFF; mem['h2B16]=8'hFF; mem['h2B17]=8'hFF;
    mem['h2B18]=8'hFF; mem['h2B19]=8'hFF; mem['h2B1A]=8'hFF; mem['h2B1B]=8'hFF;
    mem['h2B1C]=8'hFF; mem['h2B1D]=8'hFF; mem['h2B1E]=8'hFF; mem['h2B1F]=8'hFF;
    mem['h2B20]=8'hFF; mem['h2B21]=8'hFF; mem['h2B22]=8'hFF; mem['h2B23]=8'hFF;
    mem['h2B24]=8'hFF; mem['h2B25]=8'hFF; mem['h2B26]=8'hFF; mem['h2B27]=8'hFF;
    mem['h2B28]=8'hFF; mem['h2B29]=8'hFF; mem['h2B2A]=8'hFF; mem['h2B2B]=8'hFF;
    mem['h2B2C]=8'hFF; mem['h2B2D]=8'hFF; mem['h2B2E]=8'hFF; mem['h2B2F]=8'hFF;
    mem['h2B30]=8'hFF; mem['h2B31]=8'hFF; mem['h2B32]=8'hFF; mem['h2B33]=8'hFF;
    mem['h2B34]=8'hFF; mem['h2B35]=8'hFF; mem['h2B36]=8'hFF; mem['h2B37]=8'hFF;
    mem['h2B38]=8'hFF; mem['h2B39]=8'hFF; mem['h2B3A]=8'hFF; mem['h2B3B]=8'hFF;
    mem['h2B3C]=8'hFF; mem['h2B3D]=8'hFF; mem['h2B3E]=8'hFF; mem['h2B3F]=8'hFF;
    mem['h2B40]=8'hFF; mem['h2B41]=8'hFF; mem['h2B42]=8'hFF; mem['h2B43]=8'hFF;
    mem['h2B44]=8'hFF; mem['h2B45]=8'hFF; mem['h2B46]=8'hFF; mem['h2B47]=8'hFF;
    mem['h2B48]=8'hFF; mem['h2B49]=8'hFF; mem['h2B4A]=8'hFF; mem['h2B4B]=8'hFF;
    mem['h2B4C]=8'hFF; mem['h2B4D]=8'hFF; mem['h2B4E]=8'hFF; mem['h2B4F]=8'hFF;
    mem['h2B50]=8'hFF; mem['h2B51]=8'hFF; mem['h2B52]=8'hFF; mem['h2B53]=8'hFF;
    mem['h2B54]=8'hFF; mem['h2B55]=8'hFF; mem['h2B56]=8'hFF; mem['h2B57]=8'hFF;
    mem['h2B58]=8'hFF; mem['h2B59]=8'hFF; mem['h2B5A]=8'hFF; mem['h2B5B]=8'hFF;
    mem['h2B5C]=8'hFF; mem['h2B5D]=8'hFF; mem['h2B5E]=8'hFF; mem['h2B5F]=8'hFF;
    mem['h2B60]=8'hFF; mem['h2B61]=8'hFF; mem['h2B62]=8'hFF; mem['h2B63]=8'hFF;
    mem['h2B64]=8'hFF; mem['h2B65]=8'hFF; mem['h2B66]=8'hFF; mem['h2B67]=8'hFF;
    mem['h2B68]=8'hFF; mem['h2B69]=8'hFF; mem['h2B6A]=8'hFF; mem['h2B6B]=8'hFF;
    mem['h2B6C]=8'hFF; mem['h2B6D]=8'hFF; mem['h2B6E]=8'hFF; mem['h2B6F]=8'hFF;
    mem['h2B70]=8'hFF; mem['h2B71]=8'hFF; mem['h2B72]=8'hFF; mem['h2B73]=8'hFF;
    mem['h2B74]=8'hFF; mem['h2B75]=8'hFF; mem['h2B76]=8'hFF; mem['h2B77]=8'hFF;
    mem['h2B78]=8'hFF; mem['h2B79]=8'hFF; mem['h2B7A]=8'hFF; mem['h2B7B]=8'hFF;
    mem['h2B7C]=8'hFF; mem['h2B7D]=8'hFF; mem['h2B7E]=8'hFF; mem['h2B7F]=8'hFF;
    mem['h2B80]=8'hFF; mem['h2B81]=8'hFF; mem['h2B82]=8'hFF; mem['h2B83]=8'hFF;
    mem['h2B84]=8'hFF; mem['h2B85]=8'hFF; mem['h2B86]=8'hFF; mem['h2B87]=8'hFF;
    mem['h2B88]=8'hFF; mem['h2B89]=8'hFF; mem['h2B8A]=8'hFF; mem['h2B8B]=8'hFF;
    mem['h2B8C]=8'hFF; mem['h2B8D]=8'hFF; mem['h2B8E]=8'hFF; mem['h2B8F]=8'hFF;
    mem['h2B90]=8'hFF; mem['h2B91]=8'hFF; mem['h2B92]=8'hFF; mem['h2B93]=8'hFF;
    mem['h2B94]=8'hFF; mem['h2B95]=8'hFF; mem['h2B96]=8'hFF; mem['h2B97]=8'hFF;
    mem['h2B98]=8'hFF; mem['h2B99]=8'hFF; mem['h2B9A]=8'hFF; mem['h2B9B]=8'hFF;
    mem['h2B9C]=8'hFF; mem['h2B9D]=8'hFF; mem['h2B9E]=8'hFF; mem['h2B9F]=8'hFF;
    mem['h2BA0]=8'hFF; mem['h2BA1]=8'hFF; mem['h2BA2]=8'hFF; mem['h2BA3]=8'hFF;
    mem['h2BA4]=8'hFF; mem['h2BA5]=8'hFF; mem['h2BA6]=8'hFF; mem['h2BA7]=8'hFF;
    mem['h2BA8]=8'hFF; mem['h2BA9]=8'hFF; mem['h2BAA]=8'hFF; mem['h2BAB]=8'hFF;
    mem['h2BAC]=8'hFF; mem['h2BAD]=8'hFF; mem['h2BAE]=8'hFF; mem['h2BAF]=8'hFF;
    mem['h2BB0]=8'hFF; mem['h2BB1]=8'hFF; mem['h2BB2]=8'hFF; mem['h2BB3]=8'hFF;
    mem['h2BB4]=8'hFF; mem['h2BB5]=8'hFF; mem['h2BB6]=8'hFF; mem['h2BB7]=8'hFF;
    mem['h2BB8]=8'hFF; mem['h2BB9]=8'hFF; mem['h2BBA]=8'hFF; mem['h2BBB]=8'hFF;
    mem['h2BBC]=8'hFF; mem['h2BBD]=8'hFF; mem['h2BBE]=8'hFF; mem['h2BBF]=8'hFF;
    mem['h2BC0]=8'hFF; mem['h2BC1]=8'hFF; mem['h2BC2]=8'hFF; mem['h2BC3]=8'hFF;
    mem['h2BC4]=8'hFF; mem['h2BC5]=8'hFF; mem['h2BC6]=8'hFF; mem['h2BC7]=8'hFF;
    mem['h2BC8]=8'hFF; mem['h2BC9]=8'hFF; mem['h2BCA]=8'hFF; mem['h2BCB]=8'hFF;
    mem['h2BCC]=8'hFF; mem['h2BCD]=8'hFF; mem['h2BCE]=8'hFF; mem['h2BCF]=8'hFF;
    mem['h2BD0]=8'hFF; mem['h2BD1]=8'hFF; mem['h2BD2]=8'hFF; mem['h2BD3]=8'hFF;
    mem['h2BD4]=8'hFF; mem['h2BD5]=8'hFF; mem['h2BD6]=8'hFF; mem['h2BD7]=8'hFF;
    mem['h2BD8]=8'hFF; mem['h2BD9]=8'hFF; mem['h2BDA]=8'hFF; mem['h2BDB]=8'hFF;
    mem['h2BDC]=8'hFF; mem['h2BDD]=8'hFF; mem['h2BDE]=8'hFF; mem['h2BDF]=8'hFF;
    mem['h2BE0]=8'hFF; mem['h2BE1]=8'hFF; mem['h2BE2]=8'hFF; mem['h2BE3]=8'hFF;
    mem['h2BE4]=8'hFF; mem['h2BE5]=8'hFF; mem['h2BE6]=8'hFF; mem['h2BE7]=8'hFF;
    mem['h2BE8]=8'hFF; mem['h2BE9]=8'hFF; mem['h2BEA]=8'hFF; mem['h2BEB]=8'hFF;
    mem['h2BEC]=8'hFF; mem['h2BED]=8'hFF; mem['h2BEE]=8'hFF; mem['h2BEF]=8'hFF;
    mem['h2BF0]=8'hFF; mem['h2BF1]=8'hFF; mem['h2BF2]=8'hFF; mem['h2BF3]=8'hFF;
    mem['h2BF4]=8'hFF; mem['h2BF5]=8'hFF; mem['h2BF6]=8'hFF; mem['h2BF7]=8'hFF;
    mem['h2BF8]=8'hFF; mem['h2BF9]=8'hFF; mem['h2BFA]=8'hFF; mem['h2BFB]=8'hFF;
    mem['h2BFC]=8'hFF; mem['h2BFD]=8'hFF; mem['h2BFE]=8'hFF; mem['h2BFF]=8'hFF;
    mem['h2C00]=8'hFF; mem['h2C01]=8'hFF; mem['h2C02]=8'hFF; mem['h2C03]=8'hFF;
    mem['h2C04]=8'hFF; mem['h2C05]=8'hFF; mem['h2C06]=8'hFF; mem['h2C07]=8'hFF;
    mem['h2C08]=8'hFF; mem['h2C09]=8'hFF; mem['h2C0A]=8'hFF; mem['h2C0B]=8'hFF;
    mem['h2C0C]=8'hFF; mem['h2C0D]=8'hFF; mem['h2C0E]=8'hFF; mem['h2C0F]=8'hFF;
    mem['h2C10]=8'hFF; mem['h2C11]=8'hFF; mem['h2C12]=8'hFF; mem['h2C13]=8'hFF;
    mem['h2C14]=8'hFF; mem['h2C15]=8'hFF; mem['h2C16]=8'hFF; mem['h2C17]=8'hFF;
    mem['h2C18]=8'hFF; mem['h2C19]=8'hFF; mem['h2C1A]=8'hFF; mem['h2C1B]=8'hFF;
    mem['h2C1C]=8'hFF; mem['h2C1D]=8'hFF; mem['h2C1E]=8'hFF; mem['h2C1F]=8'hFF;
    mem['h2C20]=8'hFF; mem['h2C21]=8'hFF; mem['h2C22]=8'hFF; mem['h2C23]=8'hFF;
    mem['h2C24]=8'hFF; mem['h2C25]=8'hFF; mem['h2C26]=8'hFF; mem['h2C27]=8'hFF;
    mem['h2C28]=8'hFF; mem['h2C29]=8'hFF; mem['h2C2A]=8'hFF; mem['h2C2B]=8'hFF;
    mem['h2C2C]=8'hFF; mem['h2C2D]=8'hFF; mem['h2C2E]=8'hFF; mem['h2C2F]=8'hFF;
    mem['h2C30]=8'hFF; mem['h2C31]=8'hFF; mem['h2C32]=8'hFF; mem['h2C33]=8'hFF;
    mem['h2C34]=8'hFF; mem['h2C35]=8'hFF; mem['h2C36]=8'hFF; mem['h2C37]=8'hFF;
    mem['h2C38]=8'hFF; mem['h2C39]=8'hFF; mem['h2C3A]=8'hFF; mem['h2C3B]=8'hFF;
    mem['h2C3C]=8'hFF; mem['h2C3D]=8'hFF; mem['h2C3E]=8'hFF; mem['h2C3F]=8'hFF;
    mem['h2C40]=8'hFF; mem['h2C41]=8'hFF; mem['h2C42]=8'hFF; mem['h2C43]=8'hFF;
    mem['h2C44]=8'hFF; mem['h2C45]=8'hFF; mem['h2C46]=8'hFF; mem['h2C47]=8'hFF;
    mem['h2C48]=8'hFF; mem['h2C49]=8'hFF; mem['h2C4A]=8'hFF; mem['h2C4B]=8'hFF;
    mem['h2C4C]=8'hFF; mem['h2C4D]=8'hFF; mem['h2C4E]=8'hFF; mem['h2C4F]=8'hFF;
    mem['h2C50]=8'hFF; mem['h2C51]=8'hFF; mem['h2C52]=8'hFF; mem['h2C53]=8'hFF;
    mem['h2C54]=8'hFF; mem['h2C55]=8'hFF; mem['h2C56]=8'hFF; mem['h2C57]=8'hFF;
    mem['h2C58]=8'hFF; mem['h2C59]=8'hFF; mem['h2C5A]=8'hFF; mem['h2C5B]=8'hFF;
    mem['h2C5C]=8'hFF; mem['h2C5D]=8'hFF; mem['h2C5E]=8'hFF; mem['h2C5F]=8'hFF;
    mem['h2C60]=8'hFF; mem['h2C61]=8'hFF; mem['h2C62]=8'hFF; mem['h2C63]=8'hFF;
    mem['h2C64]=8'hFF; mem['h2C65]=8'hFF; mem['h2C66]=8'hFF; mem['h2C67]=8'hFF;
    mem['h2C68]=8'hFF; mem['h2C69]=8'hFF; mem['h2C6A]=8'hFF; mem['h2C6B]=8'hFF;
    mem['h2C6C]=8'hFF; mem['h2C6D]=8'hFF; mem['h2C6E]=8'hFF; mem['h2C6F]=8'hFF;
    mem['h2C70]=8'hFF; mem['h2C71]=8'hFF; mem['h2C72]=8'hFF; mem['h2C73]=8'hFF;
    mem['h2C74]=8'hFF; mem['h2C75]=8'hFF; mem['h2C76]=8'hFF; mem['h2C77]=8'hFF;
    mem['h2C78]=8'hFF; mem['h2C79]=8'hFF; mem['h2C7A]=8'hFF; mem['h2C7B]=8'hFF;
    mem['h2C7C]=8'hFF; mem['h2C7D]=8'hFF; mem['h2C7E]=8'hFF; mem['h2C7F]=8'hFF;
    mem['h2C80]=8'hFF; mem['h2C81]=8'hFF; mem['h2C82]=8'hFF; mem['h2C83]=8'hFF;
    mem['h2C84]=8'hFF; mem['h2C85]=8'hFF; mem['h2C86]=8'hFF; mem['h2C87]=8'hFF;
    mem['h2C88]=8'hFF; mem['h2C89]=8'hFF; mem['h2C8A]=8'hFF; mem['h2C8B]=8'hFF;
    mem['h2C8C]=8'hFF; mem['h2C8D]=8'hFF; mem['h2C8E]=8'hFF; mem['h2C8F]=8'hFF;
    mem['h2C90]=8'hFF; mem['h2C91]=8'hFF; mem['h2C92]=8'hFF; mem['h2C93]=8'hFF;
    mem['h2C94]=8'hFF; mem['h2C95]=8'hFF; mem['h2C96]=8'hFF; mem['h2C97]=8'hFF;
    mem['h2C98]=8'hFF; mem['h2C99]=8'hFF; mem['h2C9A]=8'hFF; mem['h2C9B]=8'hFF;
    mem['h2C9C]=8'hFF; mem['h2C9D]=8'hFF; mem['h2C9E]=8'hFF; mem['h2C9F]=8'hFF;
    mem['h2CA0]=8'hFF; mem['h2CA1]=8'hFF; mem['h2CA2]=8'hFF; mem['h2CA3]=8'hFF;
    mem['h2CA4]=8'hFF; mem['h2CA5]=8'hFF; mem['h2CA6]=8'hFF; mem['h2CA7]=8'hFF;
    mem['h2CA8]=8'hFF; mem['h2CA9]=8'hFF; mem['h2CAA]=8'hFF; mem['h2CAB]=8'hFF;
    mem['h2CAC]=8'hFF; mem['h2CAD]=8'hFF; mem['h2CAE]=8'hFF; mem['h2CAF]=8'hFF;
    mem['h2CB0]=8'hFF; mem['h2CB1]=8'hFF; mem['h2CB2]=8'hFF; mem['h2CB3]=8'hFF;
    mem['h2CB4]=8'hFF; mem['h2CB5]=8'hFF; mem['h2CB6]=8'hFF; mem['h2CB7]=8'hFF;
    mem['h2CB8]=8'hFF; mem['h2CB9]=8'hFF; mem['h2CBA]=8'hFF; mem['h2CBB]=8'hFF;
    mem['h2CBC]=8'hFF; mem['h2CBD]=8'hFF; mem['h2CBE]=8'hFF; mem['h2CBF]=8'hFF;
    mem['h2CC0]=8'hFF; mem['h2CC1]=8'hFF; mem['h2CC2]=8'hFF; mem['h2CC3]=8'hFF;
    mem['h2CC4]=8'hFF; mem['h2CC5]=8'hFF; mem['h2CC6]=8'hFF; mem['h2CC7]=8'hFF;
    mem['h2CC8]=8'hFF; mem['h2CC9]=8'hFF; mem['h2CCA]=8'hFF; mem['h2CCB]=8'hFF;
    mem['h2CCC]=8'hFF; mem['h2CCD]=8'hFF; mem['h2CCE]=8'hFF; mem['h2CCF]=8'hFF;
    mem['h2CD0]=8'hFF; mem['h2CD1]=8'hFF; mem['h2CD2]=8'hFF; mem['h2CD3]=8'hFF;
    mem['h2CD4]=8'hFF; mem['h2CD5]=8'hFF; mem['h2CD6]=8'hFF; mem['h2CD7]=8'hFF;
    mem['h2CD8]=8'hFF; mem['h2CD9]=8'hFF; mem['h2CDA]=8'hFF; mem['h2CDB]=8'hFF;
    mem['h2CDC]=8'hFF; mem['h2CDD]=8'hFF; mem['h2CDE]=8'hFF; mem['h2CDF]=8'hFF;
    mem['h2CE0]=8'hFF; mem['h2CE1]=8'hFF; mem['h2CE2]=8'hFF; mem['h2CE3]=8'hFF;
    mem['h2CE4]=8'hFF; mem['h2CE5]=8'hFF; mem['h2CE6]=8'hFF; mem['h2CE7]=8'hFF;
    mem['h2CE8]=8'hFF; mem['h2CE9]=8'hFF; mem['h2CEA]=8'hFF; mem['h2CEB]=8'hFF;
    mem['h2CEC]=8'hFF; mem['h2CED]=8'hFF; mem['h2CEE]=8'hFF; mem['h2CEF]=8'hFF;
    mem['h2CF0]=8'hFF; mem['h2CF1]=8'hFF; mem['h2CF2]=8'hFF; mem['h2CF3]=8'hFF;
    mem['h2CF4]=8'hFF; mem['h2CF5]=8'hFF; mem['h2CF6]=8'hFF; mem['h2CF7]=8'hFF;
    mem['h2CF8]=8'hFF; mem['h2CF9]=8'hFF; mem['h2CFA]=8'hFF; mem['h2CFB]=8'hFF;
    mem['h2CFC]=8'hFF; mem['h2CFD]=8'hFF; mem['h2CFE]=8'hFF; mem['h2CFF]=8'hFF;
    mem['h2D00]=8'h36; mem['h2D01]=8'h56; mem['h2D02]=8'h2E; mem['h2D03]=8'h01;
    mem['h2D04]=8'hC7; mem['h2D05]=8'hA0; mem['h2D06]=8'h70; mem['h2D07]=8'h5E;
    mem['h2D08]=8'h2D; mem['h2D09]=8'h46; mem['h2D0A]=8'h00; mem['h2D0B]=8'h10;
    mem['h2D0C]=8'h36; mem['h2D0D]=8'h54; mem['h2D0E]=8'hC7; mem['h2D0F]=8'h14;
    mem['h2D10]=8'h01; mem['h2D11]=8'h02; mem['h2D12]=8'h02; mem['h2D13]=8'hD0;
    mem['h2D14]=8'h36; mem['h2D15]=8'h83; mem['h2D16]=8'h2E; mem['h2D17]=8'h17;
    mem['h2D18]=8'hC7; mem['h2D19]=8'h2C; mem['h2D1A]=8'hFF; mem['h2D1B]=8'h02;
    mem['h2D1C]=8'h02; mem['h2D1D]=8'h04; mem['h2D1E]=8'h50; mem['h2D1F]=8'h2E;
    mem['h2D20]=8'h17; mem['h2D21]=8'hF0; mem['h2D22]=8'h30; mem['h2D23]=8'h30;
    mem['h2D24]=8'hC7; mem['h2D25]=8'h82; mem['h2D26]=8'hF0; mem['h2D27]=8'h2E;
    mem['h2D28]=8'h2F; mem['h2D29]=8'h44; mem['h2D2A]=8'hA4; mem['h2D2B]=8'h12;
    mem['h2D2C]=8'h36; mem['h2D2D]=8'h82; mem['h2D2E]=8'h2E; mem['h2D2F]=8'h17;
    mem['h2D30]=8'hCF; mem['h2D31]=8'h08; mem['h2D32]=8'hF9; mem['h2D33]=8'h16;
    mem['h2D34]=8'h02; mem['h2D35]=8'h36; mem['h2D36]=8'h4C; mem['h2D37]=8'h2E;
    mem['h2D38]=8'h17; mem['h2D39]=8'h46; mem['h2D3A]=8'h98; mem['h2D3B]=8'h07;
    mem['h2D3C]=8'h1E; mem['h2D3D]=8'h16; mem['h2D3E]=8'h26; mem['h2D3F]=8'h50;
    mem['h2D40]=8'h46; mem['h2D41]=8'hDA; mem['h2D42]=8'h02; mem['h2D43]=8'h68;
    mem['h2D44]=8'h54; mem['h2D45]=8'h2D; mem['h2D46]=8'h36; mem['h2D47]=8'h82;
    mem['h2D48]=8'h2E; mem['h2D49]=8'h17; mem['h2D4A]=8'hC7; mem['h2D4B]=8'h36;
    mem['h2D4C]=8'h3D; mem['h2D4D]=8'hBF; mem['h2D4E]=8'h48; mem['h2D4F]=8'h2C;
    mem['h2D50]=8'h2D; mem['h2D51]=8'h44; mem['h2D52]=8'h7A; mem['h2D53]=8'h07;
    mem['h2D54]=8'h36; mem['h2D55]=8'h82; mem['h2D56]=8'h2E; mem['h2D57]=8'h17;
    mem['h2D58]=8'hA8; mem['h2D59]=8'h9F; mem['h2D5A]=8'hF8; mem['h2D5B]=8'h44;
    mem['h2D5C]=8'h87; mem['h2D5D]=8'h07; mem['h2D5E]=8'h06; mem['h2D5F]=8'hCF;
    mem['h2D60]=8'h16; mem['h2D61]=8'hD2; mem['h2D62]=8'h44; mem['h2D63]=8'h96;
    mem['h2D64]=8'h02; mem['h2D65]=8'h46; mem['h2D66]=8'hAA; mem['h2D67]=8'h08;
    mem['h2D68]=8'h44; mem['h2D69]=8'h70; mem['h2D6A]=8'h2D; mem['h2D6B]=8'h36;
    mem['h2D6C]=8'h82; mem['h2D6D]=8'h44; mem['h2D6E]=8'h72; mem['h2D6F]=8'h2D;
    mem['h2D70]=8'h36; mem['h2D71]=8'h83; mem['h2D72]=8'h2E; mem['h2D73]=8'h16;
    mem['h2D74]=8'hCF; mem['h2D75]=8'h08; mem['h2D76]=8'h36; mem['h2D77]=8'hBE;
    mem['h2D78]=8'hF9; mem['h2D79]=8'h36; mem['h2D7A]=8'h86; mem['h2D7B]=8'hF9;
    mem['h2D7C]=8'h36; mem['h2D7D]=8'h86; mem['h2D7E]=8'h46; mem['h2D7F]=8'hA0;
    mem['h2D80]=8'h02; mem['h2D81]=8'h3C; mem['h2D82]=8'hA9; mem['h2D83]=8'h68;
    mem['h2D84]=8'h95; mem['h2D85]=8'h2D; mem['h2D86]=8'h36; mem['h2D87]=8'h86;
    mem['h2D88]=8'h46; mem['h2D89]=8'h03; mem['h2D8A]=8'h03; mem['h2D8B]=8'h48;
    mem['h2D8C]=8'h7C; mem['h2D8D]=8'h2D; mem['h2D8E]=8'h06; mem['h2D8F]=8'hC1;
    mem['h2D90]=8'h16; mem['h2D91]=8'hC6; mem['h2D92]=8'h44; mem['h2D93]=8'h96;
    mem['h2D94]=8'h02; mem['h2D95]=8'h36; mem['h2D96]=8'h86; mem['h2D97]=8'hCF;
    mem['h2D98]=8'h09; mem['h2D99]=8'h36; mem['h2D9A]=8'hBF; mem['h2D9B]=8'hF9;
    mem['h2D9C]=8'h36; mem['h2D9D]=8'h87; mem['h2D9E]=8'h3E; mem['h2D9F]=8'h00;
    mem['h2DA0]=8'h36; mem['h2DA1]=8'h87; mem['h2DA2]=8'h2E; mem['h2DA3]=8'h16;
    mem['h2DA4]=8'hCF; mem['h2DA5]=8'h08; mem['h2DA6]=8'hF9; mem['h2DA7]=8'h16;
    mem['h2DA8]=8'h02; mem['h2DA9]=8'h36; mem['h2DAA]=8'h4C; mem['h2DAB]=8'h2E;
    mem['h2DAC]=8'h17; mem['h2DAD]=8'h46; mem['h2DAE]=8'h98; mem['h2DAF]=8'h07;
    mem['h2DB0]=8'h26; mem['h2DB1]=8'h50; mem['h2DB2]=8'h1E; mem['h2DB3]=8'h16;
    mem['h2DB4]=8'h46; mem['h2DB5]=8'hDA; mem['h2DB6]=8'h02; mem['h2DB7]=8'h68;
    mem['h2DB8]=8'hCA; mem['h2DB9]=8'h2D; mem['h2DBA]=8'h36; mem['h2DBB]=8'h87;
    mem['h2DBC]=8'h2E; mem['h2DBD]=8'h16; mem['h2DBE]=8'hC7; mem['h2DBF]=8'h36;
    mem['h2DC0]=8'h3D; mem['h2DC1]=8'h2E; mem['h2DC2]=8'h17; mem['h2DC3]=8'hBF;
    mem['h2DC4]=8'h48; mem['h2DC5]=8'hA0; mem['h2DC6]=8'h2D; mem['h2DC7]=8'h44;
    mem['h2DC8]=8'h7A; mem['h2DC9]=8'h07; mem['h2DCA]=8'h46; mem['h2DCB]=8'h94;
    mem['h2DCC]=8'h03; mem['h2DCD]=8'h46; mem['h2DCE]=8'h00; mem['h2DCF]=8'h10;
    mem['h2DD0]=8'h36; mem['h2DD1]=8'h87; mem['h2DD2]=8'h2E; mem['h2DD3]=8'h16;
    mem['h2DD4]=8'hCF; mem['h2DD5]=8'h16; mem['h2DD6]=8'h02; mem['h2DD7]=8'h36;
    mem['h2DD8]=8'h4C; mem['h2DD9]=8'h2E; mem['h2DDA]=8'h17; mem['h2DDB]=8'h46;
    mem['h2DDC]=8'h98; mem['h2DDD]=8'h07; mem['h2DDE]=8'h30; mem['h2DDF]=8'h30;
    mem['h2DE0]=8'hD7; mem['h2DE1]=8'h36; mem['h2DE2]=8'h54; mem['h2DE3]=8'h2E;
    mem['h2DE4]=8'h01; mem['h2DE5]=8'hC7; mem['h2DE6]=8'h14; mem['h2DE7]=8'h01;
    mem['h2DE8]=8'h02; mem['h2DE9]=8'h02; mem['h2DEA]=8'h82; mem['h2DEB]=8'h36;
    mem['h2DEC]=8'h84; mem['h2DED]=8'h2E; mem['h2DEE]=8'h17; mem['h2DEF]=8'hF8;
    mem['h2DF0]=8'h36; mem['h2DF1]=8'h81; mem['h2DF2]=8'h3E; mem['h2DF3]=8'hFF;
    mem['h2DF4]=8'h07; mem['h2DF5]=8'h46; mem['h2DF6]=8'hAD; mem['h2DF7]=8'h02;
    mem['h2DF8]=8'h36; mem['h2DF9]=8'h82; mem['h2DFA]=8'hCF; mem['h2DFB]=8'h08;
    mem['h2DFC]=8'h36; mem['h2DFD]=8'h83; mem['h2DFE]=8'hF9; mem['h2DFF]=8'h36;
    mem['h2E00]=8'h83; mem['h2E01]=8'h46; mem['h2E02]=8'hA0; mem['h2E03]=8'h02;
    mem['h2E04]=8'h68; mem['h2E05]=8'h0F; mem['h2E06]=8'h2E; mem['h2E07]=8'h3C;
    mem['h2E08]=8'hA8; mem['h2E09]=8'h68; mem['h2E0A]=8'h1A; mem['h2E0B]=8'h2E;
    mem['h2E0C]=8'h46; mem['h2E0D]=8'hC8; mem['h2E0E]=8'h02; mem['h2E0F]=8'h36;
    mem['h2E10]=8'h83; mem['h2E11]=8'h46; mem['h2E12]=8'h03; mem['h2E13]=8'h03;
    mem['h2E14]=8'h48; mem['h2E15]=8'hFF; mem['h2E16]=8'h2D; mem['h2E17]=8'h44;
    mem['h2E18]=8'hDF; mem['h2E19]=8'h2E; mem['h2E1A]=8'h36; mem['h2E1B]=8'h86;
    mem['h2E1C]=8'h3E; mem['h2E1D]=8'h00; mem['h2E1E]=8'h36; mem['h2E1F]=8'h86;
    mem['h2E20]=8'h2E; mem['h2E21]=8'h16; mem['h2E22]=8'hC7; mem['h2E23]=8'h02;
    mem['h2E24]=8'h02; mem['h2E25]=8'h04; mem['h2E26]=8'h4C; mem['h2E27]=8'h2E;
    mem['h2E28]=8'h17; mem['h2E29]=8'hF0; mem['h2E2A]=8'h26; mem['h2E2B]=8'h50;
    mem['h2E2C]=8'h1E; mem['h2E2D]=8'h16; mem['h2E2E]=8'h46; mem['h2E2F]=8'hDA;
    mem['h2E30]=8'h02; mem['h2E31]=8'h68; mem['h2E32]=8'hC1; mem['h2E33]=8'h2E;
    mem['h2E34]=8'h36; mem['h2E35]=8'h86; mem['h2E36]=8'h2E; mem['h2E37]=8'h16;
    mem['h2E38]=8'hCF; mem['h2E39]=8'h08; mem['h2E3A]=8'hF9; mem['h2E3B]=8'h36;
    mem['h2E3C]=8'h3D; mem['h2E3D]=8'h2E; mem['h2E3E]=8'h17; mem['h2E3F]=8'hC7;
    mem['h2E40]=8'h09; mem['h2E41]=8'hB9; mem['h2E42]=8'h48; mem['h2E43]=8'h1E;
    mem['h2E44]=8'h2E; mem['h2E45]=8'h36; mem['h2E46]=8'h3D; mem['h2E47]=8'h2E;
    mem['h2E48]=8'h17; mem['h2E49]=8'hCF; mem['h2E4A]=8'h08; mem['h2E4B]=8'hF9;
    mem['h2E4C]=8'h36; mem['h2E4D]=8'h3E; mem['h2E4E]=8'hF9; mem['h2E4F]=8'h36;
    mem['h2E50]=8'h86; mem['h2E51]=8'h2E; mem['h2E52]=8'h16; mem['h2E53]=8'hF9;
    mem['h2E54]=8'hC7; mem['h2E55]=8'h02; mem['h2E56]=8'h02; mem['h2E57]=8'h04;
    mem['h2E58]=8'h4C; mem['h2E59]=8'hE0; mem['h2E5A]=8'h1E; mem['h2E5B]=8'h17;
    mem['h2E5C]=8'h36; mem['h2E5D]=8'h50; mem['h2E5E]=8'h2E; mem['h2E5F]=8'h16;
    mem['h2E60]=8'h46; mem['h2E61]=8'h26; mem['h2E62]=8'h0A; mem['h2E63]=8'h46;
    mem['h2E64]=8'hAD; mem['h2E65]=8'h02; mem['h2E66]=8'h36; mem['h2E67]=8'h83;
    mem['h2E68]=8'h2E; mem['h2E69]=8'h16; mem['h2E6A]=8'hCF; mem['h2E6B]=8'h08;
    mem['h2E6C]=8'h36; mem['h2E6D]=8'h84; mem['h2E6E]=8'hF9; mem['h2E6F]=8'h36;
    mem['h2E70]=8'h84; mem['h2E71]=8'h46; mem['h2E72]=8'hA0; mem['h2E73]=8'h02;
    mem['h2E74]=8'h68; mem['h2E75]=8'h89; mem['h2E76]=8'h2E; mem['h2E77]=8'h3C;
    mem['h2E78]=8'hA9; mem['h2E79]=8'h68; mem['h2E7A]=8'h94; mem['h2E7B]=8'h2E;
    mem['h2E7C]=8'h3C; mem['h2E7D]=8'hB0; mem['h2E7E]=8'h70; mem['h2E7F]=8'hDF;
    mem['h2E80]=8'h2E; mem['h2E81]=8'h3C; mem['h2E82]=8'hBA; mem['h2E83]=8'h50;
    mem['h2E84]=8'hDF; mem['h2E85]=8'h2E; mem['h2E86]=8'h46; mem['h2E87]=8'hC8;
    mem['h2E88]=8'h02; mem['h2E89]=8'h36; mem['h2E8A]=8'h84; mem['h2E8B]=8'h46;
    mem['h2E8C]=8'h03; mem['h2E8D]=8'h03; mem['h2E8E]=8'h48; mem['h2E8F]=8'h6F;
    mem['h2E90]=8'h2E; mem['h2E91]=8'h44; mem['h2E92]=8'hDF; mem['h2E93]=8'h2E;
    mem['h2E94]=8'h36; mem['h2E95]=8'h50; mem['h2E96]=8'h2E; mem['h2E97]=8'h16;
    mem['h2E98]=8'h46; mem['h2E99]=8'h24; mem['h2E9A]=8'h13; mem['h2E9B]=8'h46;
    mem['h2E9C]=8'h00; mem['h2E9D]=8'h10; mem['h2E9E]=8'h36; mem['h2E9F]=8'h54;
    mem['h2EA0]=8'hC7; mem['h2EA1]=8'h02; mem['h2EA2]=8'h02; mem['h2EA3]=8'hD0;
    mem['h2EA4]=8'h36; mem['h2EA5]=8'h3E; mem['h2EA6]=8'h2E; mem['h2EA7]=8'h17;
    mem['h2EA8]=8'hC7; mem['h2EA9]=8'h14; mem['h2EAA]=8'h01; mem['h2EAB]=8'h02;
    mem['h2EAC]=8'h02; mem['h2EAD]=8'h04; mem['h2EAE]=8'h52; mem['h2EAF]=8'hF0;
    mem['h2EB0]=8'h2E; mem['h2EB1]=8'h17; mem['h2EB2]=8'hCF; mem['h2EB3]=8'h04;
    mem['h2EB4]=8'h04; mem['h2EB5]=8'hF0; mem['h2EB6]=8'hC1; mem['h2EB7]=8'h82;
    mem['h2EB8]=8'hF8; mem['h2EB9]=8'h36; mem['h2EBA]=8'h84; mem['h2EBB]=8'h2E;
    mem['h2EBC]=8'h16; mem['h2EBD]=8'hCF; mem['h2EBE]=8'h36; mem['h2EBF]=8'h83;
    mem['h2EC0]=8'hF9; mem['h2EC1]=8'h36; mem['h2EC2]=8'h83; mem['h2EC3]=8'h46;
    mem['h2EC4]=8'hA0; mem['h2EC5]=8'h02; mem['h2EC6]=8'h3C; mem['h2EC7]=8'hAC;
    mem['h2EC8]=8'h68; mem['h2EC9]=8'hD6; mem['h2ECA]=8'h2E; mem['h2ECB]=8'h36;
    mem['h2ECC]=8'h83; mem['h2ECD]=8'h46; mem['h2ECE]=8'h03; mem['h2ECF]=8'h03;
    mem['h2ED0]=8'h48; mem['h2ED1]=8'hC1; mem['h2ED2]=8'h2E; mem['h2ED3]=8'h44;
    mem['h2ED4]=8'h4E; mem['h2ED5]=8'h0B; mem['h2ED6]=8'h36; mem['h2ED7]=8'h83;
    mem['h2ED8]=8'hCF; mem['h2ED9]=8'h36; mem['h2EDA]=8'h82; mem['h2EDB]=8'hF9;
    mem['h2EDC]=8'h44; mem['h2EDD]=8'hF5; mem['h2EDE]=8'h2D; mem['h2EDF]=8'h06;
    mem['h2EE0]=8'hC4; mem['h2EE1]=8'h16; mem['h2EE2]=8'hC5; mem['h2EE3]=8'h44;
    mem['h2EE4]=8'h96; mem['h2EE5]=8'h02; mem['h2EE6]=8'h00; mem['h2EE7]=8'h00;
end
