// rom.v
// to be included from the top module at the comple

initial
begin
    rom['h0000]=8'hC3; rom['h0001]=8'h80; rom['h0002]=8'h00; rom['h0003]=8'hFF;
    rom['h0004]=8'hFF; rom['h0005]=8'hFF; rom['h0006]=8'hFF; rom['h0007]=8'hFF;
    rom['h0008]=8'hFF; rom['h0009]=8'hFF; rom['h000A]=8'hFF; rom['h000B]=8'hFF;
    rom['h000C]=8'hFF; rom['h000D]=8'hFF; rom['h000E]=8'hFF; rom['h000F]=8'hFF;
    rom['h0010]=8'hFF; rom['h0011]=8'hFF; rom['h0012]=8'hFF; rom['h0013]=8'hFF;
    rom['h0014]=8'hFF; rom['h0015]=8'hFF; rom['h0016]=8'hFF; rom['h0017]=8'hFF;
    rom['h0018]=8'hFF; rom['h0019]=8'hFF; rom['h001A]=8'hFF; rom['h001B]=8'hFF;
    rom['h001C]=8'hFF; rom['h001D]=8'hFF; rom['h001E]=8'hFF; rom['h001F]=8'hFF;
    rom['h0020]=8'hFF; rom['h0021]=8'hFF; rom['h0022]=8'hFF; rom['h0023]=8'hFF;
    rom['h0024]=8'hFF; rom['h0025]=8'hFF; rom['h0026]=8'hFF; rom['h0027]=8'hFF;
    rom['h0028]=8'hFF; rom['h0029]=8'hFF; rom['h002A]=8'hFF; rom['h002B]=8'hFF;
    rom['h002C]=8'hFF; rom['h002D]=8'hFF; rom['h002E]=8'hFF; rom['h002F]=8'hFF;
    rom['h0030]=8'hFF; rom['h0031]=8'hFF; rom['h0032]=8'hFF; rom['h0033]=8'hFF;
    rom['h0034]=8'hFF; rom['h0035]=8'hFF; rom['h0036]=8'hFF; rom['h0037]=8'hFF;
    rom['h0038]=8'hFF; rom['h0039]=8'hFF; rom['h003A]=8'hFF; rom['h003B]=8'hFF;
    rom['h003C]=8'hFF; rom['h003D]=8'hFF; rom['h003E]=8'hFF; rom['h003F]=8'hFF;
    rom['h0040]=8'hFF; rom['h0041]=8'hFF; rom['h0042]=8'hFF; rom['h0043]=8'hFF;
    rom['h0044]=8'hFF; rom['h0045]=8'hFF; rom['h0046]=8'hFF; rom['h0047]=8'hFF;
    rom['h0048]=8'hFF; rom['h0049]=8'hFF; rom['h004A]=8'hFF; rom['h004B]=8'hFF;
    rom['h004C]=8'hFF; rom['h004D]=8'hFF; rom['h004E]=8'hFF; rom['h004F]=8'hFF;
    rom['h0050]=8'hFF; rom['h0051]=8'hFF; rom['h0052]=8'hFF; rom['h0053]=8'hFF;
    rom['h0054]=8'hFF; rom['h0055]=8'hFF; rom['h0056]=8'hFF; rom['h0057]=8'hFF;
    rom['h0058]=8'hFF; rom['h0059]=8'hFF; rom['h005A]=8'hFF; rom['h005B]=8'hFF;
    rom['h005C]=8'hFF; rom['h005D]=8'hFF; rom['h005E]=8'hFF; rom['h005F]=8'hFF;
    rom['h0060]=8'hFF; rom['h0061]=8'hFF; rom['h0062]=8'hFF; rom['h0063]=8'hFF;
    rom['h0064]=8'hFF; rom['h0065]=8'hFF; rom['h0066]=8'hFF; rom['h0067]=8'hFF;
    rom['h0068]=8'hFF; rom['h0069]=8'hFF; rom['h006A]=8'hFF; rom['h006B]=8'hFF;
    rom['h006C]=8'hFF; rom['h006D]=8'hFF; rom['h006E]=8'hFF; rom['h006F]=8'hFF;
    rom['h0070]=8'hFF; rom['h0071]=8'hFF; rom['h0072]=8'hFF; rom['h0073]=8'hFF;
    rom['h0074]=8'hFF; rom['h0075]=8'hFF; rom['h0076]=8'hFF; rom['h0077]=8'hFF;
    rom['h0078]=8'hFF; rom['h0079]=8'hFF; rom['h007A]=8'hFF; rom['h007B]=8'hFF;
    rom['h007C]=8'hFF; rom['h007D]=8'hFF; rom['h007E]=8'hFF; rom['h007F]=8'hFF;
    rom['h0080]=8'hED; rom['h0081]=8'h46; rom['h0082]=8'hF3; rom['h0083]=8'h01;
    rom['h0084]=8'h01; rom['h0085]=8'h00; rom['h0086]=8'h21; rom['h0087]=8'h00;
    rom['h0088]=8'h00; rom['h0089]=8'hAF; rom['h008A]=8'hD3; rom['h008B]=8'h0A;
    rom['h008C]=8'h78; rom['h008D]=8'hD3; rom['h008E]=8'h0B; rom['h008F]=8'h79;
    rom['h0090]=8'hD3; rom['h0091]=8'h0C; rom['h0092]=8'h7D; rom['h0093]=8'hD3;
    rom['h0094]=8'h0F; rom['h0095]=8'h7C; rom['h0096]=8'hD3; rom['h0097]=8'h10;
    rom['h0098]=8'hAF; rom['h0099]=8'hD3; rom['h009A]=8'h0D; rom['h009B]=8'hC3;
    rom['h009C]=8'h00; rom['h009D]=8'h00; rom['h009E]=8'h00; rom['h009F]=8'h00;
end
