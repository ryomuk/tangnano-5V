// rom.v
// to be included from the top module at the comple

initial
begin
    mem['h0000]=8'hF3; mem['h0001]=8'h31; mem['h0002]=8'hED; mem['h0003]=8'h80;
    mem['h0004]=8'hC3; mem['h0005]=8'h1B; mem['h0006]=8'h00; mem['h0007]=8'hFF;
    mem['h0008]=8'hC3; mem['h0009]=8'hC9; mem['h000A]=8'h00; mem['h000B]=8'hFF;
    mem['h000C]=8'hFF; mem['h000D]=8'hFF; mem['h000E]=8'hFF; mem['h000F]=8'hFF;
    mem['h0010]=8'hC3; mem['h0011]=8'h9D; mem['h0012]=8'h00; mem['h0013]=8'hFF;
    mem['h0014]=8'hFF; mem['h0015]=8'hFF; mem['h0016]=8'hFF; mem['h0017]=8'hFF;
    mem['h0018]=8'hC3; mem['h0019]=8'hC3; mem['h001A]=8'h00; mem['h001B]=8'h21;
    mem['h001C]=8'h00; mem['h001D]=8'h80; mem['h001E]=8'h11; mem['h001F]=8'h00;
    mem['h0020]=8'h80; mem['h0021]=8'h01; mem['h0022]=8'h00; mem['h0023]=8'h40;
    mem['h0024]=8'hED; mem['h0025]=8'hB0; mem['h0026]=8'hAF; mem['h0027]=8'h32;
    mem['h0028]=8'h00; mem['h0029]=8'h80; mem['h002A]=8'h32; mem['h002B]=8'h01;
    mem['h002C]=8'h80; mem['h002D]=8'h32; mem['h002E]=8'h02; mem['h002F]=8'h80;
    mem['h0030]=8'hED; mem['h0031]=8'h5E; mem['h0032]=8'h21; mem['h0033]=8'h60;
    mem['h0034]=8'h00; mem['h0035]=8'h7C; mem['h0036]=8'hED; mem['h0037]=8'h47;
    mem['h0038]=8'h21; mem['h0039]=8'h4E; mem['h003A]=8'h00; mem['h003B]=8'h0E;
    mem['h003C]=8'h01; mem['h003D]=8'h06; mem['h003E]=8'h09; mem['h003F]=8'hED;
    mem['h0040]=8'hB3; mem['h0041]=8'h21; mem['h0042]=8'h57; mem['h0043]=8'h00;
    mem['h0044]=8'h0E; mem['h0045]=8'h03; mem['h0046]=8'h06; mem['h0047]=8'h05;
    mem['h0048]=8'hED; mem['h0049]=8'hB3; mem['h004A]=8'hFB; mem['h004B]=8'hC3;
    mem['h004C]=8'hD4; mem['h004D]=8'h00; mem['h004E]=8'h18; mem['h004F]=8'h01;
    mem['h0050]=8'h14; mem['h0051]=8'h04; mem['h0052]=8'h44; mem['h0053]=8'h05;
    mem['h0054]=8'hEA; mem['h0055]=8'h03; mem['h0056]=8'hC1; mem['h0057]=8'h18;
    mem['h0058]=8'h01; mem['h0059]=8'h04; mem['h005A]=8'h02; mem['h005B]=8'h60;
    mem['h005C]=8'hFF; mem['h005D]=8'hFF; mem['h005E]=8'hFF; mem['h005F]=8'hFF;
    mem['h0060]=8'h00; mem['h0061]=8'h00; mem['h0062]=8'h00; mem['h0063]=8'h00;
    mem['h0064]=8'h00; mem['h0065]=8'h00; mem['h0066]=8'h00; mem['h0067]=8'h00;
    mem['h0068]=8'h70; mem['h0069]=8'h00; mem['h006A]=8'h70; mem['h006B]=8'h00;
    mem['h006C]=8'h73; mem['h006D]=8'h00; mem['h006E]=8'h70; mem['h006F]=8'h00;
    mem['h0070]=8'hFB; mem['h0071]=8'hED; mem['h0072]=8'h4D; mem['h0073]=8'hF5;
    mem['h0074]=8'hC5; mem['h0075]=8'hD5; mem['h0076]=8'hE5; mem['h0077]=8'hDB;
    mem['h0078]=8'h00; mem['h0079]=8'h57; mem['h007A]=8'h3A; mem['h007B]=8'h00;
    mem['h007C]=8'h80; mem['h007D]=8'hFE; mem['h007E]=8'h40; mem['h007F]=8'h28;
    mem['h0080]=8'h15; mem['h0081]=8'h3C; mem['h0082]=8'h32; mem['h0083]=8'h00;
    mem['h0084]=8'h80; mem['h0085]=8'h3A; mem['h0086]=8'h02; mem['h0087]=8'h80;
    mem['h0088]=8'h4F; mem['h0089]=8'h06; mem['h008A]=8'h00; mem['h008B]=8'h21;
    mem['h008C]=8'h03; mem['h008D]=8'h80; mem['h008E]=8'h09; mem['h008F]=8'h72;
    mem['h0090]=8'h3C; mem['h0091]=8'hE6; mem['h0092]=8'h3F; mem['h0093]=8'h32;
    mem['h0094]=8'h02; mem['h0095]=8'h80; mem['h0096]=8'hE1; mem['h0097]=8'hD1;
    mem['h0098]=8'hC1; mem['h0099]=8'hF1; mem['h009A]=8'hFB; mem['h009B]=8'hED;
    mem['h009C]=8'h4D; mem['h009D]=8'hC5; mem['h009E]=8'hD5; mem['h009F]=8'hE5;
    mem['h00A0]=8'h3A; mem['h00A1]=8'h00; mem['h00A2]=8'h80; mem['h00A3]=8'hFE;
    mem['h00A4]=8'h00; mem['h00A5]=8'h28; mem['h00A6]=8'hF9; mem['h00A7]=8'hF3;
    mem['h00A8]=8'h3D; mem['h00A9]=8'h32; mem['h00AA]=8'h00; mem['h00AB]=8'h80;
    mem['h00AC]=8'h3A; mem['h00AD]=8'h01; mem['h00AE]=8'h80; mem['h00AF]=8'h4F;
    mem['h00B0]=8'h06; mem['h00B1]=8'h00; mem['h00B2]=8'h21; mem['h00B3]=8'h03;
    mem['h00B4]=8'h80; mem['h00B5]=8'h09; mem['h00B6]=8'h56; mem['h00B7]=8'h3C;
    mem['h00B8]=8'hE6; mem['h00B9]=8'h3F; mem['h00BA]=8'h32; mem['h00BB]=8'h01;
    mem['h00BC]=8'h80; mem['h00BD]=8'h7A; mem['h00BE]=8'hFB; mem['h00BF]=8'hE1;
    mem['h00C0]=8'hD1; mem['h00C1]=8'hC1; mem['h00C2]=8'hC9; mem['h00C3]=8'h3A;
    mem['h00C4]=8'h00; mem['h00C5]=8'h80; mem['h00C6]=8'hFE; mem['h00C7]=8'h00;
    mem['h00C8]=8'hC9; mem['h00C9]=8'hF5; mem['h00CA]=8'hDB; mem['h00CB]=8'h01;
    mem['h00CC]=8'hCB; mem['h00CD]=8'h57; mem['h00CE]=8'h28; mem['h00CF]=8'hFA;
    mem['h00D0]=8'hF1; mem['h00D1]=8'hD3; mem['h00D2]=8'h00; mem['h00D3]=8'hC9;
    mem['h00D4]=8'hC3; mem['h00D5]=8'hDA; mem['h00D6]=8'h00; mem['h00D7]=8'hC3;
    mem['h00D8]=8'h4F; mem['h00D9]=8'h01; mem['h00DA]=8'hC3; mem['h00DB]=8'hE1;
    mem['h00DC]=8'h00; mem['h00DD]=8'h92; mem['h00DE]=8'h09; mem['h00DF]=8'h08;
    mem['h00E0]=8'h11; mem['h00E1]=8'h21; mem['h00E2]=8'h45; mem['h00E3]=8'h80;
    mem['h00E4]=8'hF9; mem['h00E5]=8'hC3; mem['h00E6]=8'h23; mem['h00E7]=8'h1D;
    mem['h00E8]=8'h11; mem['h00E9]=8'hB9; mem['h00EA]=8'h03; mem['h00EB]=8'h06;
    mem['h00EC]=8'h63; mem['h00ED]=8'h21; mem['h00EE]=8'h45; mem['h00EF]=8'h80;
    mem['h00F0]=8'h1A; mem['h00F1]=8'h77; mem['h00F2]=8'h23; mem['h00F3]=8'h13;
    mem['h00F4]=8'h05; mem['h00F5]=8'hC2; mem['h00F6]=8'hF0; mem['h00F7]=8'h00;
    mem['h00F8]=8'hF9; mem['h00F9]=8'hCD; mem['h00FA]=8'hBA; mem['h00FB]=8'h05;
    mem['h00FC]=8'hCD; mem['h00FD]=8'h88; mem['h00FE]=8'h0B; mem['h00FF]=8'h32;
    mem['h0100]=8'hEF; mem['h0101]=8'h80; mem['h0102]=8'h32; mem['h0103]=8'h3E;
    mem['h0104]=8'h81; mem['h0105]=8'h21; mem['h0106]=8'hA2; mem['h0107]=8'h81;
    mem['h0108]=8'h23; mem['h0109]=8'h7C; mem['h010A]=8'hB5; mem['h010B]=8'hCA;
    mem['h010C]=8'h17; mem['h010D]=8'h01; mem['h010E]=8'h7E; mem['h010F]=8'h47;
    mem['h0110]=8'h2F; mem['h0111]=8'h77; mem['h0112]=8'hBE; mem['h0113]=8'h70;
    mem['h0114]=8'hCA; mem['h0115]=8'h08; mem['h0116]=8'h01; mem['h0117]=8'h2B;
    mem['h0118]=8'h11; mem['h0119]=8'hA1; mem['h011A]=8'h81; mem['h011B]=8'hCD;
    mem['h011C]=8'h50; mem['h011D]=8'h07; mem['h011E]=8'hDA; mem['h011F]=8'h58;
    mem['h0120]=8'h01; mem['h0121]=8'h11; mem['h0122]=8'hCE; mem['h0123]=8'hFF;
    mem['h0124]=8'h22; mem['h0125]=8'hF4; mem['h0126]=8'h80; mem['h0127]=8'h19;
    mem['h0128]=8'h22; mem['h0129]=8'h9F; mem['h012A]=8'h80; mem['h012B]=8'hCD;
    mem['h012C]=8'h95; mem['h012D]=8'h05; mem['h012E]=8'h2A; mem['h012F]=8'h9F;
    mem['h0130]=8'h80; mem['h0131]=8'h11; mem['h0132]=8'hEF; mem['h0133]=8'hFF;
    mem['h0134]=8'h19; mem['h0135]=8'h11; mem['h0136]=8'h3E; mem['h0137]=8'h81;
    mem['h0138]=8'h7D; mem['h0139]=8'h93; mem['h013A]=8'h6F; mem['h013B]=8'h7C;
    mem['h013C]=8'h9A; mem['h013D]=8'h67; mem['h013E]=8'hE5; mem['h013F]=8'h21;
    mem['h0140]=8'h70; mem['h0141]=8'h01; mem['h0142]=8'hCD; mem['h0143]=8'h26;
    mem['h0144]=8'h12; mem['h0145]=8'hE1; mem['h0146]=8'hCD; mem['h0147]=8'hC9;
    mem['h0148]=8'h18; mem['h0149]=8'h21; mem['h014A]=8'h61; mem['h014B]=8'h01;
    mem['h014C]=8'hCD; mem['h014D]=8'h26; mem['h014E]=8'h12; mem['h014F]=8'h31;
    mem['h0150]=8'hAB; mem['h0151]=8'h80; mem['h0152]=8'hCD; mem['h0153]=8'hBA;
    mem['h0154]=8'h05; mem['h0155]=8'hC3; mem['h0156]=8'hD3; mem['h0157]=8'h04;
    mem['h0158]=8'h21; mem['h0159]=8'hA7; mem['h015A]=8'h01; mem['h015B]=8'hCD;
    mem['h015C]=8'h26; mem['h015D]=8'h12; mem['h015E]=8'hC3; mem['h015F]=8'h5E;
    mem['h0160]=8'h01; mem['h0161]=8'h20; mem['h0162]=8'h42; mem['h0163]=8'h79;
    mem['h0164]=8'h74; mem['h0165]=8'h65; mem['h0166]=8'h73; mem['h0167]=8'h20;
    mem['h0168]=8'h66; mem['h0169]=8'h72; mem['h016A]=8'h65; mem['h016B]=8'h65;
    mem['h016C]=8'h0D; mem['h016D]=8'h0A; mem['h016E]=8'h00; mem['h016F]=8'h00;
    mem['h0170]=8'h5A; mem['h0171]=8'h38; mem['h0172]=8'h30; mem['h0173]=8'h20;
    mem['h0174]=8'h42; mem['h0175]=8'h41; mem['h0176]=8'h53; mem['h0177]=8'h49;
    mem['h0178]=8'h43; mem['h0179]=8'h20; mem['h017A]=8'h56; mem['h017B]=8'h65;
    mem['h017C]=8'h72; mem['h017D]=8'h20; mem['h017E]=8'h34; mem['h017F]=8'h2E;
    mem['h0180]=8'h37; mem['h0181]=8'h62; mem['h0182]=8'h0D; mem['h0183]=8'h0A;
    mem['h0184]=8'h43; mem['h0185]=8'h6F; mem['h0186]=8'h70; mem['h0187]=8'h79;
    mem['h0188]=8'h72; mem['h0189]=8'h69; mem['h018A]=8'h67; mem['h018B]=8'h68;
    mem['h018C]=8'h74; mem['h018D]=8'h20; mem['h018E]=8'h28; mem['h018F]=8'h43;
    mem['h0190]=8'h29; mem['h0191]=8'h20; mem['h0192]=8'h31; mem['h0193]=8'h39;
    mem['h0194]=8'h37; mem['h0195]=8'h38; mem['h0196]=8'h20; mem['h0197]=8'h62;
    mem['h0198]=8'h79; mem['h0199]=8'h20; mem['h019A]=8'h4D; mem['h019B]=8'h69;
    mem['h019C]=8'h63; mem['h019D]=8'h72; mem['h019E]=8'h6F; mem['h019F]=8'h73;
    mem['h01A0]=8'h6F; mem['h01A1]=8'h66; mem['h01A2]=8'h74; mem['h01A3]=8'h0D;
    mem['h01A4]=8'h0A; mem['h01A5]=8'h00; mem['h01A6]=8'h00; mem['h01A7]=8'h4D;
    mem['h01A8]=8'h65; mem['h01A9]=8'h6D; mem['h01AA]=8'h6F; mem['h01AB]=8'h72;
    mem['h01AC]=8'h79; mem['h01AD]=8'h20; mem['h01AE]=8'h73; mem['h01AF]=8'h69;
    mem['h01B0]=8'h7A; mem['h01B1]=8'h65; mem['h01B2]=8'h20; mem['h01B3]=8'h6E;
    mem['h01B4]=8'h6F; mem['h01B5]=8'h74; mem['h01B6]=8'h20; mem['h01B7]=8'h65;
    mem['h01B8]=8'h6E; mem['h01B9]=8'h6F; mem['h01BA]=8'h75; mem['h01BB]=8'h67;
    mem['h01BC]=8'h68; mem['h01BD]=8'h0D; mem['h01BE]=8'h0A; mem['h01BF]=8'h54;
    mem['h01C0]=8'h68; mem['h01C1]=8'h65; mem['h01C2]=8'h20; mem['h01C3]=8'h73;
    mem['h01C4]=8'h79; mem['h01C5]=8'h73; mem['h01C6]=8'h74; mem['h01C7]=8'h65;
    mem['h01C8]=8'h6D; mem['h01C9]=8'h20; mem['h01CA]=8'h69; mem['h01CB]=8'h73;
    mem['h01CC]=8'h20; mem['h01CD]=8'h73; mem['h01CE]=8'h74; mem['h01CF]=8'h6F;
    mem['h01D0]=8'h70; mem['h01D1]=8'h70; mem['h01D2]=8'h65; mem['h01D3]=8'h64;
    mem['h01D4]=8'h2E; mem['h01D5]=8'h0D; mem['h01D6]=8'h0A; mem['h01D7]=8'h00;
    mem['h01D8]=8'h00; mem['h01D9]=8'h3E; mem['h01DA]=8'h17; mem['h01DB]=8'h02;
    mem['h01DC]=8'h18; mem['h01DD]=8'h54; mem['h01DE]=8'h17; mem['h01DF]=8'h48;
    mem['h01E0]=8'h80; mem['h01E1]=8'hE6; mem['h01E2]=8'h10; mem['h01E3]=8'h6B;
    mem['h01E4]=8'h14; mem['h01E5]=8'h14; mem['h01E6]=8'h11; mem['h01E7]=8'hC8;
    mem['h01E8]=8'h19; mem['h01E9]=8'hA7; mem['h01EA]=8'h1A; mem['h01EB]=8'hE3;
    mem['h01EC]=8'h15; mem['h01ED]=8'h16; mem['h01EE]=8'h1A; mem['h01EF]=8'h1C;
    mem['h01F0]=8'h1B; mem['h01F1]=8'h22; mem['h01F2]=8'h1B; mem['h01F3]=8'h83;
    mem['h01F4]=8'h1B; mem['h01F5]=8'h98; mem['h01F6]=8'h1B; mem['h01F7]=8'hBF;
    mem['h01F8]=8'h14; mem['h01F9]=8'h03; mem['h01FA]=8'h1C; mem['h01FB]=8'h96;
    mem['h01FC]=8'h80; mem['h01FD]=8'h98; mem['h01FE]=8'h13; mem['h01FF]=8'hB0;
    mem['h0200]=8'h11; mem['h0201]=8'h32; mem['h0202]=8'h14; mem['h0203]=8'hA7;
    mem['h0204]=8'h13; mem['h0205]=8'hB8; mem['h0206]=8'h13; mem['h0207]=8'h25;
    mem['h0208]=8'h1C; mem['h0209]=8'hB8; mem['h020A]=8'h1C; mem['h020B]=8'hC8;
    mem['h020C]=8'h13; mem['h020D]=8'hF8; mem['h020E]=8'h13; mem['h020F]=8'h02;
    mem['h0210]=8'h14; mem['h0211]=8'hC5; mem['h0212]=8'h4E; mem['h0213]=8'h44;
    mem['h0214]=8'hC6; mem['h0215]=8'h4F; mem['h0216]=8'h52; mem['h0217]=8'hCE;
    mem['h0218]=8'h45; mem['h0219]=8'h58; mem['h021A]=8'h54; mem['h021B]=8'hC4;
    mem['h021C]=8'h41; mem['h021D]=8'h54; mem['h021E]=8'h41; mem['h021F]=8'hC9;
    mem['h0220]=8'h4E; mem['h0221]=8'h50; mem['h0222]=8'h55; mem['h0223]=8'h54;
    mem['h0224]=8'hC4; mem['h0225]=8'h49; mem['h0226]=8'h4D; mem['h0227]=8'hD2;
    mem['h0228]=8'h45; mem['h0229]=8'h41; mem['h022A]=8'h44; mem['h022B]=8'hCC;
    mem['h022C]=8'h45; mem['h022D]=8'h54; mem['h022E]=8'hC7; mem['h022F]=8'h4F;
    mem['h0230]=8'h54; mem['h0231]=8'h4F; mem['h0232]=8'hD2; mem['h0233]=8'h55;
    mem['h0234]=8'h4E; mem['h0235]=8'hC9; mem['h0236]=8'h46; mem['h0237]=8'hD2;
    mem['h0238]=8'h45; mem['h0239]=8'h53; mem['h023A]=8'h54; mem['h023B]=8'h4F;
    mem['h023C]=8'h52; mem['h023D]=8'h45; mem['h023E]=8'hC7; mem['h023F]=8'h4F;
    mem['h0240]=8'h53; mem['h0241]=8'h55; mem['h0242]=8'h42; mem['h0243]=8'hD2;
    mem['h0244]=8'h45; mem['h0245]=8'h54; mem['h0246]=8'h55; mem['h0247]=8'h52;
    mem['h0248]=8'h4E; mem['h0249]=8'hD2; mem['h024A]=8'h45; mem['h024B]=8'h4D;
    mem['h024C]=8'hD3; mem['h024D]=8'h54; mem['h024E]=8'h4F; mem['h024F]=8'h50;
    mem['h0250]=8'hCF; mem['h0251]=8'h55; mem['h0252]=8'h54; mem['h0253]=8'hCF;
    mem['h0254]=8'h4E; mem['h0255]=8'hCE; mem['h0256]=8'h55; mem['h0257]=8'h4C;
    mem['h0258]=8'h4C; mem['h0259]=8'hD7; mem['h025A]=8'h41; mem['h025B]=8'h49;
    mem['h025C]=8'h54; mem['h025D]=8'hC4; mem['h025E]=8'h45; mem['h025F]=8'h46;
    mem['h0260]=8'hD0; mem['h0261]=8'h4F; mem['h0262]=8'h4B; mem['h0263]=8'h45;
    mem['h0264]=8'hC4; mem['h0265]=8'h4F; mem['h0266]=8'h4B; mem['h0267]=8'h45;
    mem['h0268]=8'hD3; mem['h0269]=8'h43; mem['h026A]=8'h52; mem['h026B]=8'h45;
    mem['h026C]=8'h45; mem['h026D]=8'h4E; mem['h026E]=8'hCC; mem['h026F]=8'h49;
    mem['h0270]=8'h4E; mem['h0271]=8'h45; mem['h0272]=8'h53; mem['h0273]=8'hC3;
    mem['h0274]=8'h4C; mem['h0275]=8'h53; mem['h0276]=8'hD7; mem['h0277]=8'h49;
    mem['h0278]=8'h44; mem['h0279]=8'h54; mem['h027A]=8'h48; mem['h027B]=8'hCD;
    mem['h027C]=8'h4F; mem['h027D]=8'h4E; mem['h027E]=8'h49; mem['h027F]=8'h54;
    mem['h0280]=8'h4F; mem['h0281]=8'h52; mem['h0282]=8'hD3; mem['h0283]=8'h45;
    mem['h0284]=8'h54; mem['h0285]=8'hD2; mem['h0286]=8'h45; mem['h0287]=8'h53;
    mem['h0288]=8'h45; mem['h0289]=8'h54; mem['h028A]=8'hD0; mem['h028B]=8'h52;
    mem['h028C]=8'h49; mem['h028D]=8'h4E; mem['h028E]=8'h54; mem['h028F]=8'hC3;
    mem['h0290]=8'h4F; mem['h0291]=8'h4E; mem['h0292]=8'h54; mem['h0293]=8'hCC;
    mem['h0294]=8'h49; mem['h0295]=8'h53; mem['h0296]=8'h54; mem['h0297]=8'hC3;
    mem['h0298]=8'h4C; mem['h0299]=8'h45; mem['h029A]=8'h41; mem['h029B]=8'h52;
    mem['h029C]=8'hC3; mem['h029D]=8'h4C; mem['h029E]=8'h4F; mem['h029F]=8'h41;
    mem['h02A0]=8'h44; mem['h02A1]=8'hC3; mem['h02A2]=8'h53; mem['h02A3]=8'h41;
    mem['h02A4]=8'h56; mem['h02A5]=8'h45; mem['h02A6]=8'hCE; mem['h02A7]=8'h45;
    mem['h02A8]=8'h57; mem['h02A9]=8'hD4; mem['h02AA]=8'h41; mem['h02AB]=8'h42;
    mem['h02AC]=8'h28; mem['h02AD]=8'hD4; mem['h02AE]=8'h4F; mem['h02AF]=8'hC6;
    mem['h02B0]=8'h4E; mem['h02B1]=8'hD3; mem['h02B2]=8'h50; mem['h02B3]=8'h43;
    mem['h02B4]=8'h28; mem['h02B5]=8'hD4; mem['h02B6]=8'h48; mem['h02B7]=8'h45;
    mem['h02B8]=8'h4E; mem['h02B9]=8'hCE; mem['h02BA]=8'h4F; mem['h02BB]=8'h54;
    mem['h02BC]=8'hD3; mem['h02BD]=8'h54; mem['h02BE]=8'h45; mem['h02BF]=8'h50;
    mem['h02C0]=8'hAB; mem['h02C1]=8'hAD; mem['h02C2]=8'hAA; mem['h02C3]=8'hAF;
    mem['h02C4]=8'hDE; mem['h02C5]=8'hC1; mem['h02C6]=8'h4E; mem['h02C7]=8'h44;
    mem['h02C8]=8'hCF; mem['h02C9]=8'h52; mem['h02CA]=8'hBE; mem['h02CB]=8'hBD;
    mem['h02CC]=8'hBC; mem['h02CD]=8'hD3; mem['h02CE]=8'h47; mem['h02CF]=8'h4E;
    mem['h02D0]=8'hC9; mem['h02D1]=8'h4E; mem['h02D2]=8'h54; mem['h02D3]=8'hC1;
    mem['h02D4]=8'h42; mem['h02D5]=8'h53; mem['h02D6]=8'hD5; mem['h02D7]=8'h53;
    mem['h02D8]=8'h52; mem['h02D9]=8'hC6; mem['h02DA]=8'h52; mem['h02DB]=8'h45;
    mem['h02DC]=8'hC9; mem['h02DD]=8'h4E; mem['h02DE]=8'h50; mem['h02DF]=8'hD0;
    mem['h02E0]=8'h4F; mem['h02E1]=8'h53; mem['h02E2]=8'hD3; mem['h02E3]=8'h51;
    mem['h02E4]=8'h52; mem['h02E5]=8'hD2; mem['h02E6]=8'h4E; mem['h02E7]=8'h44;
    mem['h02E8]=8'hCC; mem['h02E9]=8'h4F; mem['h02EA]=8'h47; mem['h02EB]=8'hC5;
    mem['h02EC]=8'h58; mem['h02ED]=8'h50; mem['h02EE]=8'hC3; mem['h02EF]=8'h4F;
    mem['h02F0]=8'h53; mem['h02F1]=8'hD3; mem['h02F2]=8'h49; mem['h02F3]=8'h4E;
    mem['h02F4]=8'hD4; mem['h02F5]=8'h41; mem['h02F6]=8'h4E; mem['h02F7]=8'hC1;
    mem['h02F8]=8'h54; mem['h02F9]=8'h4E; mem['h02FA]=8'hD0; mem['h02FB]=8'h45;
    mem['h02FC]=8'h45; mem['h02FD]=8'h4B; mem['h02FE]=8'hC4; mem['h02FF]=8'h45;
    mem['h0300]=8'h45; mem['h0301]=8'h4B; mem['h0302]=8'hD0; mem['h0303]=8'h4F;
    mem['h0304]=8'h49; mem['h0305]=8'h4E; mem['h0306]=8'h54; mem['h0307]=8'hCC;
    mem['h0308]=8'h45; mem['h0309]=8'h4E; mem['h030A]=8'hD3; mem['h030B]=8'h54;
    mem['h030C]=8'h52; mem['h030D]=8'h24; mem['h030E]=8'hD6; mem['h030F]=8'h41;
    mem['h0310]=8'h4C; mem['h0311]=8'hC1; mem['h0312]=8'h53; mem['h0313]=8'h43;
    mem['h0314]=8'hC3; mem['h0315]=8'h48; mem['h0316]=8'h52; mem['h0317]=8'h24;
    mem['h0318]=8'hC8; mem['h0319]=8'h45; mem['h031A]=8'h58; mem['h031B]=8'h24;
    mem['h031C]=8'hC2; mem['h031D]=8'h49; mem['h031E]=8'h4E; mem['h031F]=8'h24;
    mem['h0320]=8'hCC; mem['h0321]=8'h45; mem['h0322]=8'h46; mem['h0323]=8'h54;
    mem['h0324]=8'h24; mem['h0325]=8'hD2; mem['h0326]=8'h49; mem['h0327]=8'h47;
    mem['h0328]=8'h48; mem['h0329]=8'h54; mem['h032A]=8'h24; mem['h032B]=8'hCD;
    mem['h032C]=8'h49; mem['h032D]=8'h44; mem['h032E]=8'h24; mem['h032F]=8'h80;
    mem['h0330]=8'h2A; mem['h0331]=8'h09; mem['h0332]=8'h27; mem['h0333]=8'h08;
    mem['h0334]=8'h02; mem['h0335]=8'h0D; mem['h0336]=8'h77; mem['h0337]=8'h0A;
    mem['h0338]=8'h09; mem['h0339]=8'h0C; mem['h033A]=8'h3E; mem['h033B]=8'h0F;
    mem['h033C]=8'h38; mem['h033D]=8'h0C; mem['h033E]=8'h8E; mem['h033F]=8'h0A;
    mem['h0340]=8'h34; mem['h0341]=8'h0A; mem['h0342]=8'h17; mem['h0343]=8'h0A;
    mem['h0344]=8'h06; mem['h0345]=8'h0B; mem['h0346]=8'hF0; mem['h0347]=8'h08;
    mem['h0348]=8'h23; mem['h0349]=8'h0A; mem['h034A]=8'h52; mem['h034B]=8'h0A;
    mem['h034C]=8'h79; mem['h034D]=8'h0A; mem['h034E]=8'h28; mem['h034F]=8'h09;
    mem['h0350]=8'h77; mem['h0351]=8'h14; mem['h0352]=8'hE8; mem['h0353]=8'h0A;
    mem['h0354]=8'h69; mem['h0355]=8'h09; mem['h0356]=8'h7D; mem['h0357]=8'h14;
    mem['h0358]=8'h1C; mem['h0359]=8'h11; mem['h035A]=8'hC6; mem['h035B]=8'h14;
    mem['h035C]=8'h0E; mem['h035D]=8'h1C; mem['h035E]=8'h79; mem['h035F]=8'h0A;
    mem['h0360]=8'hF4; mem['h0361]=8'h1B; mem['h0362]=8'hE7; mem['h0363]=8'h1B;
    mem['h0364]=8'hEC; mem['h0365]=8'h1B; mem['h0366]=8'h20; mem['h0367]=8'h1D;
    mem['h0368]=8'h99; mem['h0369]=8'h80; mem['h036A]=8'h9C; mem['h036B]=8'h80;
    mem['h036C]=8'h2A; mem['h036D]=8'h0B; mem['h036E]=8'h56; mem['h036F]=8'h09;
    mem['h0370]=8'h9C; mem['h0371]=8'h07; mem['h0372]=8'hD1; mem['h0373]=8'h09;
    mem['h0374]=8'h79; mem['h0375]=8'h0A; mem['h0376]=8'h79; mem['h0377]=8'h0A;
    mem['h0378]=8'h94; mem['h0379]=8'h05; mem['h037A]=8'h79; mem['h037B]=8'hB0;
    mem['h037C]=8'h18; mem['h037D]=8'h79; mem['h037E]=8'hE4; mem['h037F]=8'h14;
    mem['h0380]=8'h7C; mem['h0381]=8'h22; mem['h0382]=8'h16; mem['h0383]=8'h7C;
    mem['h0384]=8'h83; mem['h0385]=8'h16; mem['h0386]=8'h7F; mem['h0387]=8'hD1;
    mem['h0388]=8'h19; mem['h0389]=8'h50; mem['h038A]=8'h97; mem['h038B]=8'h0E;
    mem['h038C]=8'h46; mem['h038D]=8'h96; mem['h038E]=8'h0E; mem['h038F]=8'h4E;
    mem['h0390]=8'h46; mem['h0391]=8'h53; mem['h0392]=8'h4E; mem['h0393]=8'h52;
    mem['h0394]=8'h47; mem['h0395]=8'h4F; mem['h0396]=8'h44; mem['h0397]=8'h46;
    mem['h0398]=8'h43; mem['h0399]=8'h4F; mem['h039A]=8'h56; mem['h039B]=8'h4F;
    mem['h039C]=8'h4D; mem['h039D]=8'h55; mem['h039E]=8'h4C; mem['h039F]=8'h42;
    mem['h03A0]=8'h53; mem['h03A1]=8'h44; mem['h03A2]=8'h44; mem['h03A3]=8'h2F;
    mem['h03A4]=8'h30; mem['h03A5]=8'h49; mem['h03A6]=8'h44; mem['h03A7]=8'h54;
    mem['h03A8]=8'h4D; mem['h03A9]=8'h4F; mem['h03AA]=8'h53; mem['h03AB]=8'h4C;
    mem['h03AC]=8'h53; mem['h03AD]=8'h53; mem['h03AE]=8'h54; mem['h03AF]=8'h43;
    mem['h03B0]=8'h4E; mem['h03B1]=8'h55; mem['h03B2]=8'h46; mem['h03B3]=8'h4D;
    mem['h03B4]=8'h4F; mem['h03B5]=8'h48; mem['h03B6]=8'h58; mem['h03B7]=8'h42;
    mem['h03B8]=8'h4E; mem['h03B9]=8'hC3; mem['h03BA]=8'h4F; mem['h03BB]=8'h01;
    mem['h03BC]=8'hC3; mem['h03BD]=8'hA7; mem['h03BE]=8'h09; mem['h03BF]=8'hD3;
    mem['h03C0]=8'h00; mem['h03C1]=8'hC9; mem['h03C2]=8'hD6; mem['h03C3]=8'h00;
    mem['h03C4]=8'h6F; mem['h03C5]=8'h7C; mem['h03C6]=8'hDE; mem['h03C7]=8'h00;
    mem['h03C8]=8'h67; mem['h03C9]=8'h78; mem['h03CA]=8'hDE; mem['h03CB]=8'h00;
    mem['h03CC]=8'h47; mem['h03CD]=8'h3E; mem['h03CE]=8'h00; mem['h03CF]=8'hC9;
    mem['h03D0]=8'h00; mem['h03D1]=8'h00; mem['h03D2]=8'h00; mem['h03D3]=8'h35;
    mem['h03D4]=8'h4A; mem['h03D5]=8'hCA; mem['h03D6]=8'h99; mem['h03D7]=8'h39;
    mem['h03D8]=8'h1C; mem['h03D9]=8'h76; mem['h03DA]=8'h98; mem['h03DB]=8'h22;
    mem['h03DC]=8'h95; mem['h03DD]=8'hB3; mem['h03DE]=8'h98; mem['h03DF]=8'h0A;
    mem['h03E0]=8'hDD; mem['h03E1]=8'h47; mem['h03E2]=8'h98; mem['h03E3]=8'h53;
    mem['h03E4]=8'hD1; mem['h03E5]=8'h99; mem['h03E6]=8'h99; mem['h03E7]=8'h0A;
    mem['h03E8]=8'h1A; mem['h03E9]=8'h9F; mem['h03EA]=8'h98; mem['h03EB]=8'h65;
    mem['h03EC]=8'hBC; mem['h03ED]=8'hCD; mem['h03EE]=8'h98; mem['h03EF]=8'hD6;
    mem['h03F0]=8'h77; mem['h03F1]=8'h3E; mem['h03F2]=8'h98; mem['h03F3]=8'h52;
    mem['h03F4]=8'hC7; mem['h03F5]=8'h4F; mem['h03F6]=8'h80; mem['h03F7]=8'hDB;
    mem['h03F8]=8'h00; mem['h03F9]=8'hC9; mem['h03FA]=8'h01; mem['h03FB]=8'hFF;
    mem['h03FC]=8'h1C; mem['h03FD]=8'h00; mem['h03FE]=8'h00; mem['h03FF]=8'h14;
    mem['h0400]=8'h00; mem['h0401]=8'h14; mem['h0402]=8'h00; mem['h0403]=8'h00;
    mem['h0404]=8'h00; mem['h0405]=8'h00; mem['h0406]=8'h00; mem['h0407]=8'hC3;
    mem['h0408]=8'hCD; mem['h0409]=8'h06; mem['h040A]=8'hC3; mem['h040B]=8'h00;
    mem['h040C]=8'h00; mem['h040D]=8'hC3; mem['h040E]=8'h00; mem['h040F]=8'h00;
    mem['h0410]=8'hC3; mem['h0411]=8'h00; mem['h0412]=8'h00; mem['h0413]=8'hA2;
    mem['h0414]=8'h81; mem['h0415]=8'hFE; mem['h0416]=8'hFF; mem['h0417]=8'h3F;
    mem['h0418]=8'h81; mem['h0419]=8'h20; mem['h041A]=8'h45; mem['h041B]=8'h72;
    mem['h041C]=8'h72; mem['h041D]=8'h6F; mem['h041E]=8'h72; mem['h041F]=8'h00;
    mem['h0420]=8'h20; mem['h0421]=8'h69; mem['h0422]=8'h6E; mem['h0423]=8'h20;
    mem['h0424]=8'h00; mem['h0425]=8'h4F; mem['h0426]=8'h6B; mem['h0427]=8'h0D;
    mem['h0428]=8'h0A; mem['h0429]=8'h00; mem['h042A]=8'h00; mem['h042B]=8'h42;
    mem['h042C]=8'h72; mem['h042D]=8'h65; mem['h042E]=8'h61; mem['h042F]=8'h6B;
    mem['h0430]=8'h00; mem['h0431]=8'h21; mem['h0432]=8'h04; mem['h0433]=8'h00;
    mem['h0434]=8'h39; mem['h0435]=8'h7E; mem['h0436]=8'h23; mem['h0437]=8'hFE;
    mem['h0438]=8'h81; mem['h0439]=8'hC0; mem['h043A]=8'h4E; mem['h043B]=8'h23;
    mem['h043C]=8'h46; mem['h043D]=8'h23; mem['h043E]=8'hE5; mem['h043F]=8'h69;
    mem['h0440]=8'h60; mem['h0441]=8'h7A; mem['h0442]=8'hB3; mem['h0443]=8'hEB;
    mem['h0444]=8'hCA; mem['h0445]=8'h4B; mem['h0446]=8'h04; mem['h0447]=8'hEB;
    mem['h0448]=8'hCD; mem['h0449]=8'h50; mem['h044A]=8'h07; mem['h044B]=8'h01;
    mem['h044C]=8'h0D; mem['h044D]=8'h00; mem['h044E]=8'hE1; mem['h044F]=8'hC8;
    mem['h0450]=8'h09; mem['h0451]=8'hC3; mem['h0452]=8'h35; mem['h0453]=8'h04;
    mem['h0454]=8'hCD; mem['h0455]=8'h6E; mem['h0456]=8'h04; mem['h0457]=8'hC5;
    mem['h0458]=8'hE3; mem['h0459]=8'hC1; mem['h045A]=8'hCD; mem['h045B]=8'h50;
    mem['h045C]=8'h07; mem['h045D]=8'h7E; mem['h045E]=8'h02; mem['h045F]=8'hC8;
    mem['h0460]=8'h0B; mem['h0461]=8'h2B; mem['h0462]=8'hC3; mem['h0463]=8'h5A;
    mem['h0464]=8'h04; mem['h0465]=8'hE5; mem['h0466]=8'h2A; mem['h0467]=8'h1F;
    mem['h0468]=8'h81; mem['h0469]=8'h06; mem['h046A]=8'h00; mem['h046B]=8'h09;
    mem['h046C]=8'h09; mem['h046D]=8'h3E; mem['h046E]=8'hE5; mem['h046F]=8'h3E;
    mem['h0470]=8'hD0; mem['h0471]=8'h95; mem['h0472]=8'h6F; mem['h0473]=8'h3E;
    mem['h0474]=8'hFF; mem['h0475]=8'h9C; mem['h0476]=8'hDA; mem['h0477]=8'h7D;
    mem['h0478]=8'h04; mem['h0479]=8'h67; mem['h047A]=8'h39; mem['h047B]=8'hE1;
    mem['h047C]=8'hD8; mem['h047D]=8'h1E; mem['h047E]=8'h0C; mem['h047F]=8'hC3;
    mem['h0480]=8'h9C; mem['h0481]=8'h04; mem['h0482]=8'h2A; mem['h0483]=8'h0E;
    mem['h0484]=8'h81; mem['h0485]=8'h22; mem['h0486]=8'hA1; mem['h0487]=8'h80;
    mem['h0488]=8'h1E; mem['h0489]=8'h02; mem['h048A]=8'h01; mem['h048B]=8'h1E;
    mem['h048C]=8'h14; mem['h048D]=8'h01; mem['h048E]=8'h1E; mem['h048F]=8'h00;
    mem['h0490]=8'h01; mem['h0491]=8'h1E; mem['h0492]=8'h12; mem['h0493]=8'h01;
    mem['h0494]=8'h1E; mem['h0495]=8'h22; mem['h0496]=8'h01; mem['h0497]=8'h1E;
    mem['h0498]=8'h0A; mem['h0499]=8'h01; mem['h049A]=8'h1E; mem['h049B]=8'h18;
    mem['h049C]=8'hCD; mem['h049D]=8'hBA; mem['h049E]=8'h05; mem['h049F]=8'h32;
    mem['h04A0]=8'h8A; mem['h04A1]=8'h80; mem['h04A2]=8'hCD; mem['h04A3]=8'h7B;
    mem['h04A4]=8'h0B; mem['h04A5]=8'h21; mem['h04A6]=8'h8F; mem['h04A7]=8'h03;
    mem['h04A8]=8'h57; mem['h04A9]=8'h3E; mem['h04AA]=8'h3F; mem['h04AB]=8'hCD;
    mem['h04AC]=8'h61; mem['h04AD]=8'h07; mem['h04AE]=8'h19; mem['h04AF]=8'h7E;
    mem['h04B0]=8'hCD; mem['h04B1]=8'h61; mem['h04B2]=8'h07; mem['h04B3]=8'hCD;
    mem['h04B4]=8'hE0; mem['h04B5]=8'h08; mem['h04B6]=8'hCD; mem['h04B7]=8'h61;
    mem['h04B8]=8'h07; mem['h04B9]=8'h21; mem['h04BA]=8'h19; mem['h04BB]=8'h04;
    mem['h04BC]=8'hCD; mem['h04BD]=8'h26; mem['h04BE]=8'h12; mem['h04BF]=8'h2A;
    mem['h04C0]=8'hA1; mem['h04C1]=8'h80; mem['h04C2]=8'h11; mem['h04C3]=8'hFE;
    mem['h04C4]=8'hFF; mem['h04C5]=8'hCD; mem['h04C6]=8'h50; mem['h04C7]=8'h07;
    mem['h04C8]=8'hCA; mem['h04C9]=8'hE1; mem['h04CA]=8'h00; mem['h04CB]=8'h7C;
    mem['h04CC]=8'hA5; mem['h04CD]=8'h3C; mem['h04CE]=8'hC4; mem['h04CF]=8'hC1;
    mem['h04D0]=8'h18; mem['h04D1]=8'h3E; mem['h04D2]=8'hC1; mem['h04D3]=8'hAF;
    mem['h04D4]=8'h32; mem['h04D5]=8'h8A; mem['h04D6]=8'h80; mem['h04D7]=8'hCD;
    mem['h04D8]=8'h7B; mem['h04D9]=8'h0B; mem['h04DA]=8'h21; mem['h04DB]=8'h25;
    mem['h04DC]=8'h04; mem['h04DD]=8'hCD; mem['h04DE]=8'h26; mem['h04DF]=8'h12;
    mem['h04E0]=8'h21; mem['h04E1]=8'hFF; mem['h04E2]=8'hFF; mem['h04E3]=8'h22;
    mem['h04E4]=8'hA1; mem['h04E5]=8'h80; mem['h04E6]=8'hCD; mem['h04E7]=8'hCD;
    mem['h04E8]=8'h06; mem['h04E9]=8'hDA; mem['h04EA]=8'hE0; mem['h04EB]=8'h04;
    mem['h04EC]=8'hCD; mem['h04ED]=8'hE0; mem['h04EE]=8'h08; mem['h04EF]=8'h3C;
    mem['h04F0]=8'h3D; mem['h04F1]=8'hCA; mem['h04F2]=8'hE0; mem['h04F3]=8'h04;
    mem['h04F4]=8'hF5; mem['h04F5]=8'hCD; mem['h04F6]=8'hAC; mem['h04F7]=8'h09;
    mem['h04F8]=8'hD5; mem['h04F9]=8'hCD; mem['h04FA]=8'hE4; mem['h04FB]=8'h05;
    mem['h04FC]=8'h47; mem['h04FD]=8'hD1; mem['h04FE]=8'hF1; mem['h04FF]=8'hD2;
    mem['h0500]=8'hC0; mem['h0501]=8'h08; mem['h0502]=8'hD5; mem['h0503]=8'hC5;
    mem['h0504]=8'hAF; mem['h0505]=8'h32; mem['h0506]=8'h11; mem['h0507]=8'h81;
    mem['h0508]=8'hCD; mem['h0509]=8'hE0; mem['h050A]=8'h08; mem['h050B]=8'hB7;
    mem['h050C]=8'hF5; mem['h050D]=8'hCD; mem['h050E]=8'h74; mem['h050F]=8'h05;
    mem['h0510]=8'hDA; mem['h0511]=8'h19; mem['h0512]=8'h05; mem['h0513]=8'hF1;
    mem['h0514]=8'hF5; mem['h0515]=8'hCA; mem['h0516]=8'h4D; mem['h0517]=8'h0A;
    mem['h0518]=8'hB7; mem['h0519]=8'hC5; mem['h051A]=8'hD2; mem['h051B]=8'h30;
    mem['h051C]=8'h05; mem['h051D]=8'hEB; mem['h051E]=8'h2A; mem['h051F]=8'h1B;
    mem['h0520]=8'h81; mem['h0521]=8'h1A; mem['h0522]=8'h02; mem['h0523]=8'h03;
    mem['h0524]=8'h13; mem['h0525]=8'hCD; mem['h0526]=8'h50; mem['h0527]=8'h07;
    mem['h0528]=8'hC2; mem['h0529]=8'h21; mem['h052A]=8'h05; mem['h052B]=8'h60;
    mem['h052C]=8'h69; mem['h052D]=8'h22; mem['h052E]=8'h1B; mem['h052F]=8'h81;
    mem['h0530]=8'hD1; mem['h0531]=8'hF1; mem['h0532]=8'hCA; mem['h0533]=8'h57;
    mem['h0534]=8'h05; mem['h0535]=8'h2A; mem['h0536]=8'h1B; mem['h0537]=8'h81;
    mem['h0538]=8'hE3; mem['h0539]=8'hC1; mem['h053A]=8'h09; mem['h053B]=8'hE5;
    mem['h053C]=8'hCD; mem['h053D]=8'h54; mem['h053E]=8'h04; mem['h053F]=8'hE1;
    mem['h0540]=8'h22; mem['h0541]=8'h1B; mem['h0542]=8'h81; mem['h0543]=8'hEB;
    mem['h0544]=8'h74; mem['h0545]=8'hD1; mem['h0546]=8'h23; mem['h0547]=8'h23;
    mem['h0548]=8'h73; mem['h0549]=8'h23; mem['h054A]=8'h72; mem['h054B]=8'h23;
    mem['h054C]=8'h11; mem['h054D]=8'hA6; mem['h054E]=8'h80; mem['h054F]=8'h1A;
    mem['h0550]=8'h77; mem['h0551]=8'h23; mem['h0552]=8'h13; mem['h0553]=8'hB7;
    mem['h0554]=8'hC2; mem['h0555]=8'h4F; mem['h0556]=8'h05; mem['h0557]=8'hCD;
    mem['h0558]=8'hA0; mem['h0559]=8'h05; mem['h055A]=8'h23; mem['h055B]=8'hEB;
    mem['h055C]=8'h62; mem['h055D]=8'h6B; mem['h055E]=8'h7E; mem['h055F]=8'h23;
    mem['h0560]=8'hB6; mem['h0561]=8'hCA; mem['h0562]=8'hE0; mem['h0563]=8'h04;
    mem['h0564]=8'h23; mem['h0565]=8'h23; mem['h0566]=8'h23; mem['h0567]=8'hAF;
    mem['h0568]=8'hBE; mem['h0569]=8'h23; mem['h056A]=8'hC2; mem['h056B]=8'h68;
    mem['h056C]=8'h05; mem['h056D]=8'hEB; mem['h056E]=8'h73; mem['h056F]=8'h23;
    mem['h0570]=8'h72; mem['h0571]=8'hC3; mem['h0572]=8'h5C; mem['h0573]=8'h05;
    mem['h0574]=8'h2A; mem['h0575]=8'hA3; mem['h0576]=8'h80; mem['h0577]=8'h44;
    mem['h0578]=8'h4D; mem['h0579]=8'h7E; mem['h057A]=8'h23; mem['h057B]=8'hB6;
    mem['h057C]=8'h2B; mem['h057D]=8'hC8; mem['h057E]=8'h23; mem['h057F]=8'h23;
    mem['h0580]=8'h7E; mem['h0581]=8'h23; mem['h0582]=8'h66; mem['h0583]=8'h6F;
    mem['h0584]=8'hCD; mem['h0585]=8'h50; mem['h0586]=8'h07; mem['h0587]=8'h60;
    mem['h0588]=8'h69; mem['h0589]=8'h7E; mem['h058A]=8'h23; mem['h058B]=8'h66;
    mem['h058C]=8'h6F; mem['h058D]=8'h3F; mem['h058E]=8'hC8; mem['h058F]=8'h3F;
    mem['h0590]=8'hD0; mem['h0591]=8'hC3; mem['h0592]=8'h77; mem['h0593]=8'h05;
    mem['h0594]=8'hC0; mem['h0595]=8'h2A; mem['h0596]=8'hA3; mem['h0597]=8'h80;
    mem['h0598]=8'hAF; mem['h0599]=8'h77; mem['h059A]=8'h23; mem['h059B]=8'h77;
    mem['h059C]=8'h23; mem['h059D]=8'h22; mem['h059E]=8'h1B; mem['h059F]=8'h81;
    mem['h05A0]=8'h2A; mem['h05A1]=8'hA3; mem['h05A2]=8'h80; mem['h05A3]=8'h2B;
    mem['h05A4]=8'h22; mem['h05A5]=8'h13; mem['h05A6]=8'h81; mem['h05A7]=8'h2A;
    mem['h05A8]=8'hF4; mem['h05A9]=8'h80; mem['h05AA]=8'h22; mem['h05AB]=8'h08;
    mem['h05AC]=8'h81; mem['h05AD]=8'hAF; mem['h05AE]=8'hCD; mem['h05AF]=8'hF0;
    mem['h05B0]=8'h08; mem['h05B1]=8'h2A; mem['h05B2]=8'h1B; mem['h05B3]=8'h81;
    mem['h05B4]=8'h22; mem['h05B5]=8'h1D; mem['h05B6]=8'h81; mem['h05B7]=8'h22;
    mem['h05B8]=8'h1F; mem['h05B9]=8'h81; mem['h05BA]=8'hC1; mem['h05BB]=8'h2A;
    mem['h05BC]=8'h9F; mem['h05BD]=8'h80; mem['h05BE]=8'hF9; mem['h05BF]=8'h21;
    mem['h05C0]=8'hF8; mem['h05C1]=8'h80; mem['h05C2]=8'h22; mem['h05C3]=8'hF6;
    mem['h05C4]=8'h80; mem['h05C5]=8'hAF; mem['h05C6]=8'h6F; mem['h05C7]=8'h67;
    mem['h05C8]=8'h22; mem['h05C9]=8'h19; mem['h05CA]=8'h81; mem['h05CB]=8'h32;
    mem['h05CC]=8'h10; mem['h05CD]=8'h81; mem['h05CE]=8'h22; mem['h05CF]=8'h23;
    mem['h05D0]=8'h81; mem['h05D1]=8'hE5; mem['h05D2]=8'hC5; mem['h05D3]=8'h2A;
    mem['h05D4]=8'h13; mem['h05D5]=8'h81; mem['h05D6]=8'hC9; mem['h05D7]=8'h3E;
    mem['h05D8]=8'h3F; mem['h05D9]=8'hCD; mem['h05DA]=8'h61; mem['h05DB]=8'h07;
    mem['h05DC]=8'h3E; mem['h05DD]=8'h20; mem['h05DE]=8'hCD; mem['h05DF]=8'h61;
    mem['h05E0]=8'h07; mem['h05E1]=8'hC3; mem['h05E2]=8'h93; mem['h05E3]=8'h80;
    mem['h05E4]=8'hAF; mem['h05E5]=8'h32; mem['h05E6]=8'hF3; mem['h05E7]=8'h80;
    mem['h05E8]=8'h0E; mem['h05E9]=8'h05; mem['h05EA]=8'h11; mem['h05EB]=8'hA6;
    mem['h05EC]=8'h80; mem['h05ED]=8'h7E; mem['h05EE]=8'hFE; mem['h05EF]=8'h20;
    mem['h05F0]=8'hCA; mem['h05F1]=8'h6C; mem['h05F2]=8'h06; mem['h05F3]=8'h47;
    mem['h05F4]=8'hFE; mem['h05F5]=8'h22; mem['h05F6]=8'hCA; mem['h05F7]=8'h8C;
    mem['h05F8]=8'h06; mem['h05F9]=8'hB7; mem['h05FA]=8'hCA; mem['h05FB]=8'h93;
    mem['h05FC]=8'h06; mem['h05FD]=8'h3A; mem['h05FE]=8'hF3; mem['h05FF]=8'h80;
    mem['h0600]=8'hB7; mem['h0601]=8'h7E; mem['h0602]=8'hC2; mem['h0603]=8'h6C;
    mem['h0604]=8'h06; mem['h0605]=8'hFE; mem['h0606]=8'h3F; mem['h0607]=8'h3E;
    mem['h0608]=8'h9E; mem['h0609]=8'hCA; mem['h060A]=8'h6C; mem['h060B]=8'h06;
    mem['h060C]=8'h7E; mem['h060D]=8'hFE; mem['h060E]=8'h30; mem['h060F]=8'hDA;
    mem['h0610]=8'h17; mem['h0611]=8'h06; mem['h0612]=8'hFE; mem['h0613]=8'h3C;
    mem['h0614]=8'hDA; mem['h0615]=8'h6C; mem['h0616]=8'h06; mem['h0617]=8'hD5;
    mem['h0618]=8'h11; mem['h0619]=8'h10; mem['h061A]=8'h02; mem['h061B]=8'hC5;
    mem['h061C]=8'h01; mem['h061D]=8'h68; mem['h061E]=8'h06; mem['h061F]=8'hC5;
    mem['h0620]=8'h06; mem['h0621]=8'h7F; mem['h0622]=8'h7E; mem['h0623]=8'hFE;
    mem['h0624]=8'h61; mem['h0625]=8'hDA; mem['h0626]=8'h30; mem['h0627]=8'h06;
    mem['h0628]=8'hFE; mem['h0629]=8'h7B; mem['h062A]=8'hD2; mem['h062B]=8'h30;
    mem['h062C]=8'h06; mem['h062D]=8'hE6; mem['h062E]=8'h5F; mem['h062F]=8'h77;
    mem['h0630]=8'h4E; mem['h0631]=8'hEB; mem['h0632]=8'h23; mem['h0633]=8'hB6;
    mem['h0634]=8'hF2; mem['h0635]=8'h32; mem['h0636]=8'h06; mem['h0637]=8'h04;
    mem['h0638]=8'h7E; mem['h0639]=8'hE6; mem['h063A]=8'h7F; mem['h063B]=8'hC8;
    mem['h063C]=8'hB9; mem['h063D]=8'hC2; mem['h063E]=8'h32; mem['h063F]=8'h06;
    mem['h0640]=8'hEB; mem['h0641]=8'hE5; mem['h0642]=8'h13; mem['h0643]=8'h1A;
    mem['h0644]=8'hB7; mem['h0645]=8'hFA; mem['h0646]=8'h64; mem['h0647]=8'h06;
    mem['h0648]=8'h4F; mem['h0649]=8'h78; mem['h064A]=8'hFE; mem['h064B]=8'h88;
    mem['h064C]=8'hC2; mem['h064D]=8'h53; mem['h064E]=8'h06; mem['h064F]=8'hCD;
    mem['h0650]=8'hE0; mem['h0651]=8'h08; mem['h0652]=8'h2B; mem['h0653]=8'h23;
    mem['h0654]=8'h7E; mem['h0655]=8'hFE; mem['h0656]=8'h61; mem['h0657]=8'hDA;
    mem['h0658]=8'h5C; mem['h0659]=8'h06; mem['h065A]=8'hE6; mem['h065B]=8'h5F;
    mem['h065C]=8'hB9; mem['h065D]=8'hCA; mem['h065E]=8'h42; mem['h065F]=8'h06;
    mem['h0660]=8'hE1; mem['h0661]=8'hC3; mem['h0662]=8'h30; mem['h0663]=8'h06;
    mem['h0664]=8'h48; mem['h0665]=8'hF1; mem['h0666]=8'hEB; mem['h0667]=8'hC9;
    mem['h0668]=8'hEB; mem['h0669]=8'h79; mem['h066A]=8'hC1; mem['h066B]=8'hD1;
    mem['h066C]=8'h23; mem['h066D]=8'h12; mem['h066E]=8'h13; mem['h066F]=8'h0C;
    mem['h0670]=8'hD6; mem['h0671]=8'h3A; mem['h0672]=8'hCA; mem['h0673]=8'h7A;
    mem['h0674]=8'h06; mem['h0675]=8'hFE; mem['h0676]=8'h49; mem['h0677]=8'hC2;
    mem['h0678]=8'h7D; mem['h0679]=8'h06; mem['h067A]=8'h32; mem['h067B]=8'hF3;
    mem['h067C]=8'h80; mem['h067D]=8'hD6; mem['h067E]=8'h54; mem['h067F]=8'hC2;
    mem['h0680]=8'hED; mem['h0681]=8'h05; mem['h0682]=8'h47; mem['h0683]=8'h7E;
    mem['h0684]=8'hB7; mem['h0685]=8'hCA; mem['h0686]=8'h93; mem['h0687]=8'h06;
    mem['h0688]=8'hB8; mem['h0689]=8'hCA; mem['h068A]=8'h6C; mem['h068B]=8'h06;
    mem['h068C]=8'h23; mem['h068D]=8'h12; mem['h068E]=8'h0C; mem['h068F]=8'h13;
    mem['h0690]=8'hC3; mem['h0691]=8'h83; mem['h0692]=8'h06; mem['h0693]=8'h21;
    mem['h0694]=8'hA5; mem['h0695]=8'h80; mem['h0696]=8'h12; mem['h0697]=8'h13;
    mem['h0698]=8'h12; mem['h0699]=8'h13; mem['h069A]=8'h12; mem['h069B]=8'hC9;
    mem['h069C]=8'h3A; mem['h069D]=8'h89; mem['h069E]=8'h80; mem['h069F]=8'hB7;
    mem['h06A0]=8'h3E; mem['h06A1]=8'h00; mem['h06A2]=8'h32; mem['h06A3]=8'h89;
    mem['h06A4]=8'h80; mem['h06A5]=8'hC2; mem['h06A6]=8'hB0; mem['h06A7]=8'h06;
    mem['h06A8]=8'h05; mem['h06A9]=8'hCA; mem['h06AA]=8'hCD; mem['h06AB]=8'h06;
    mem['h06AC]=8'hCD; mem['h06AD]=8'h61; mem['h06AE]=8'h07; mem['h06AF]=8'h3E;
    mem['h06B0]=8'h05; mem['h06B1]=8'h2B; mem['h06B2]=8'hCA; mem['h06B3]=8'hC4;
    mem['h06B4]=8'h06; mem['h06B5]=8'h7E; mem['h06B6]=8'hCD; mem['h06B7]=8'h61;
    mem['h06B8]=8'h07; mem['h06B9]=8'hC3; mem['h06BA]=8'hD6; mem['h06BB]=8'h06;
    mem['h06BC]=8'h05; mem['h06BD]=8'h2B; mem['h06BE]=8'hCD; mem['h06BF]=8'h61;
    mem['h06C0]=8'h07; mem['h06C1]=8'hC2; mem['h06C2]=8'hD6; mem['h06C3]=8'h06;
    mem['h06C4]=8'hCD; mem['h06C5]=8'h61; mem['h06C6]=8'h07; mem['h06C7]=8'hCD;
    mem['h06C8]=8'h88; mem['h06C9]=8'h0B; mem['h06CA]=8'hC3; mem['h06CB]=8'hCD;
    mem['h06CC]=8'h06; mem['h06CD]=8'h21; mem['h06CE]=8'hA6; mem['h06CF]=8'h80;
    mem['h06D0]=8'h06; mem['h06D1]=8'h01; mem['h06D2]=8'hAF; mem['h06D3]=8'h32;
    mem['h06D4]=8'h89; mem['h06D5]=8'h80; mem['h06D6]=8'hCD; mem['h06D7]=8'h8B;
    mem['h06D8]=8'h07; mem['h06D9]=8'h4F; mem['h06DA]=8'hFE; mem['h06DB]=8'h7F;
    mem['h06DC]=8'hCA; mem['h06DD]=8'h9C; mem['h06DE]=8'h06; mem['h06DF]=8'h3A;
    mem['h06E0]=8'h89; mem['h06E1]=8'h80; mem['h06E2]=8'hB7; mem['h06E3]=8'hCA;
    mem['h06E4]=8'hEF; mem['h06E5]=8'h06; mem['h06E6]=8'h3E; mem['h06E7]=8'h00;
    mem['h06E8]=8'hCD; mem['h06E9]=8'h61; mem['h06EA]=8'h07; mem['h06EB]=8'hAF;
    mem['h06EC]=8'h32; mem['h06ED]=8'h89; mem['h06EE]=8'h80; mem['h06EF]=8'h79;
    mem['h06F0]=8'hFE; mem['h06F1]=8'h07; mem['h06F2]=8'hCA; mem['h06F3]=8'h33;
    mem['h06F4]=8'h07; mem['h06F5]=8'hFE; mem['h06F6]=8'h03; mem['h06F7]=8'hCC;
    mem['h06F8]=8'h88; mem['h06F9]=8'h0B; mem['h06FA]=8'h37; mem['h06FB]=8'hC8;
    mem['h06FC]=8'hFE; mem['h06FD]=8'h0D; mem['h06FE]=8'hCA; mem['h06FF]=8'h83;
    mem['h0700]=8'h0B; mem['h0701]=8'hFE; mem['h0702]=8'h15; mem['h0703]=8'hCA;
    mem['h0704]=8'hC7; mem['h0705]=8'h06; mem['h0706]=8'hFE; mem['h0707]=8'h40;
    mem['h0708]=8'hCA; mem['h0709]=8'hC4; mem['h070A]=8'h06; mem['h070B]=8'hFE;
    mem['h070C]=8'h5F; mem['h070D]=8'hCA; mem['h070E]=8'hBC; mem['h070F]=8'h06;
    mem['h0710]=8'hFE; mem['h0711]=8'h08; mem['h0712]=8'hCA; mem['h0713]=8'hBC;
    mem['h0714]=8'h06; mem['h0715]=8'hFE; mem['h0716]=8'h12; mem['h0717]=8'hC2;
    mem['h0718]=8'h2E; mem['h0719]=8'h07; mem['h071A]=8'hC5; mem['h071B]=8'hD5;
    mem['h071C]=8'hE5; mem['h071D]=8'h36; mem['h071E]=8'h00; mem['h071F]=8'hCD;
    mem['h0720]=8'h32; mem['h0721]=8'h1D; mem['h0722]=8'h21; mem['h0723]=8'hA6;
    mem['h0724]=8'h80; mem['h0725]=8'hCD; mem['h0726]=8'h26; mem['h0727]=8'h12;
    mem['h0728]=8'hE1; mem['h0729]=8'hD1; mem['h072A]=8'hC1; mem['h072B]=8'hC3;
    mem['h072C]=8'hD6; mem['h072D]=8'h06; mem['h072E]=8'hFE; mem['h072F]=8'h20;
    mem['h0730]=8'hDA; mem['h0731]=8'hD6; mem['h0732]=8'h06; mem['h0733]=8'h78;
    mem['h0734]=8'hFE; mem['h0735]=8'h49; mem['h0736]=8'h3E; mem['h0737]=8'h07;
    mem['h0738]=8'hD2; mem['h0739]=8'h48; mem['h073A]=8'h07; mem['h073B]=8'h79;
    mem['h073C]=8'h71; mem['h073D]=8'h32; mem['h073E]=8'h11; mem['h073F]=8'h81;
    mem['h0740]=8'h23; mem['h0741]=8'h04; mem['h0742]=8'hCD; mem['h0743]=8'h61;
    mem['h0744]=8'h07; mem['h0745]=8'hC3; mem['h0746]=8'hD6; mem['h0747]=8'h06;
    mem['h0748]=8'hCD; mem['h0749]=8'h61; mem['h074A]=8'h07; mem['h074B]=8'h3E;
    mem['h074C]=8'h08; mem['h074D]=8'hC3; mem['h074E]=8'h42; mem['h074F]=8'h07;
    mem['h0750]=8'h7C; mem['h0751]=8'h92; mem['h0752]=8'hC0; mem['h0753]=8'h7D;
    mem['h0754]=8'h93; mem['h0755]=8'hC9; mem['h0756]=8'h7E; mem['h0757]=8'hE3;
    mem['h0758]=8'hBE; mem['h0759]=8'h23; mem['h075A]=8'hE3; mem['h075B]=8'hCA;
    mem['h075C]=8'hE0; mem['h075D]=8'h08; mem['h075E]=8'hC3; mem['h075F]=8'h88;
    mem['h0760]=8'h04; mem['h0761]=8'hF5; mem['h0762]=8'h3A; mem['h0763]=8'h8A;
    mem['h0764]=8'h80; mem['h0765]=8'hB7; mem['h0766]=8'hC2; mem['h0767]=8'h5B;
    mem['h0768]=8'h12; mem['h0769]=8'hF1; mem['h076A]=8'hC5; mem['h076B]=8'hF5;
    mem['h076C]=8'hFE; mem['h076D]=8'h20; mem['h076E]=8'hDA; mem['h076F]=8'h85;
    mem['h0770]=8'h07; mem['h0771]=8'h3A; mem['h0772]=8'h87; mem['h0773]=8'h80;
    mem['h0774]=8'h47; mem['h0775]=8'h3A; mem['h0776]=8'hF0; mem['h0777]=8'h80;
    mem['h0778]=8'h04; mem['h0779]=8'hCA; mem['h077A]=8'h81; mem['h077B]=8'h07;
    mem['h077C]=8'h05; mem['h077D]=8'hB8; mem['h077E]=8'hCC; mem['h077F]=8'h88;
    mem['h0780]=8'h0B; mem['h0781]=8'h3C; mem['h0782]=8'h32; mem['h0783]=8'hF0;
    mem['h0784]=8'h80; mem['h0785]=8'hF1; mem['h0786]=8'hC1; mem['h0787]=8'hCD;
    mem['h0788]=8'h1D; mem['h0789]=8'h1D; mem['h078A]=8'hC9; mem['h078B]=8'hCD;
    mem['h078C]=8'hE5; mem['h078D]=8'h1B; mem['h078E]=8'hE6; mem['h078F]=8'h7F;
    mem['h0790]=8'hFE; mem['h0791]=8'h0F; mem['h0792]=8'hC0; mem['h0793]=8'h3A;
    mem['h0794]=8'h8A; mem['h0795]=8'h80; mem['h0796]=8'h2F; mem['h0797]=8'h32;
    mem['h0798]=8'h8A; mem['h0799]=8'h80; mem['h079A]=8'hAF; mem['h079B]=8'hC9;
    mem['h079C]=8'hCD; mem['h079D]=8'hAC; mem['h079E]=8'h09; mem['h079F]=8'hC0;
    mem['h07A0]=8'hC1; mem['h07A1]=8'hCD; mem['h07A2]=8'h74; mem['h07A3]=8'h05;
    mem['h07A4]=8'hC5; mem['h07A5]=8'hCD; mem['h07A6]=8'hF2; mem['h07A7]=8'h07;
    mem['h07A8]=8'hE1; mem['h07A9]=8'h4E; mem['h07AA]=8'h23; mem['h07AB]=8'h46;
    mem['h07AC]=8'h23; mem['h07AD]=8'h78; mem['h07AE]=8'hB1; mem['h07AF]=8'hCA;
    mem['h07B0]=8'hD3; mem['h07B1]=8'h04; mem['h07B2]=8'hCD; mem['h07B3]=8'hFB;
    mem['h07B4]=8'h07; mem['h07B5]=8'hCD; mem['h07B6]=8'h0B; mem['h07B7]=8'h09;
    mem['h07B8]=8'hC5; mem['h07B9]=8'hCD; mem['h07BA]=8'h88; mem['h07BB]=8'h0B;
    mem['h07BC]=8'h5E; mem['h07BD]=8'h23; mem['h07BE]=8'h56; mem['h07BF]=8'h23;
    mem['h07C0]=8'hE5; mem['h07C1]=8'hEB; mem['h07C2]=8'hCD; mem['h07C3]=8'hC9;
    mem['h07C4]=8'h18; mem['h07C5]=8'h3E; mem['h07C6]=8'h20; mem['h07C7]=8'hE1;
    mem['h07C8]=8'hCD; mem['h07C9]=8'h61; mem['h07CA]=8'h07; mem['h07CB]=8'h7E;
    mem['h07CC]=8'hB7; mem['h07CD]=8'h23; mem['h07CE]=8'hCA; mem['h07CF]=8'hA8;
    mem['h07D0]=8'h07; mem['h07D1]=8'hF2; mem['h07D2]=8'hC8; mem['h07D3]=8'h07;
    mem['h07D4]=8'hD6; mem['h07D5]=8'h7F; mem['h07D6]=8'h4F; mem['h07D7]=8'h11;
    mem['h07D8]=8'h11; mem['h07D9]=8'h02; mem['h07DA]=8'h1A; mem['h07DB]=8'h13;
    mem['h07DC]=8'hB7; mem['h07DD]=8'hF2; mem['h07DE]=8'hDA; mem['h07DF]=8'h07;
    mem['h07E0]=8'h0D; mem['h07E1]=8'hC2; mem['h07E2]=8'hDA; mem['h07E3]=8'h07;
    mem['h07E4]=8'hE6; mem['h07E5]=8'h7F; mem['h07E6]=8'hCD; mem['h07E7]=8'h61;
    mem['h07E8]=8'h07; mem['h07E9]=8'h1A; mem['h07EA]=8'h13; mem['h07EB]=8'hB7;
    mem['h07EC]=8'hF2; mem['h07ED]=8'hE4; mem['h07EE]=8'h07; mem['h07EF]=8'hC3;
    mem['h07F0]=8'hCB; mem['h07F1]=8'h07; mem['h07F2]=8'hE5; mem['h07F3]=8'h2A;
    mem['h07F4]=8'h8D; mem['h07F5]=8'h80; mem['h07F6]=8'h22; mem['h07F7]=8'h8B;
    mem['h07F8]=8'h80; mem['h07F9]=8'hE1; mem['h07FA]=8'hC9; mem['h07FB]=8'hE5;
    mem['h07FC]=8'hD5; mem['h07FD]=8'h2A; mem['h07FE]=8'h8B; mem['h07FF]=8'h80;
    mem['h0800]=8'h11; mem['h0801]=8'hFF; mem['h0802]=8'hFF; mem['h0803]=8'hED;
    mem['h0804]=8'h5A; mem['h0805]=8'h22; mem['h0806]=8'h8B; mem['h0807]=8'h80;
    mem['h0808]=8'hD1; mem['h0809]=8'hE1; mem['h080A]=8'hF0; mem['h080B]=8'hE5;
    mem['h080C]=8'h2A; mem['h080D]=8'h8D; mem['h080E]=8'h80; mem['h080F]=8'h22;
    mem['h0810]=8'h8B; mem['h0811]=8'h80; mem['h0812]=8'hCD; mem['h0813]=8'hE5;
    mem['h0814]=8'h1B; mem['h0815]=8'hFE; mem['h0816]=8'h03; mem['h0817]=8'hCA;
    mem['h0818]=8'h1E; mem['h0819]=8'h08; mem['h081A]=8'hE1; mem['h081B]=8'hC3;
    mem['h081C]=8'hFB; mem['h081D]=8'h07; mem['h081E]=8'h2A; mem['h081F]=8'h8D;
    mem['h0820]=8'h80; mem['h0821]=8'h22; mem['h0822]=8'h8B; mem['h0823]=8'h80;
    mem['h0824]=8'hC3; mem['h0825]=8'h52; mem['h0826]=8'h01; mem['h0827]=8'h3E;
    mem['h0828]=8'h64; mem['h0829]=8'h32; mem['h082A]=8'h10; mem['h082B]=8'h81;
    mem['h082C]=8'hCD; mem['h082D]=8'h8E; mem['h082E]=8'h0A; mem['h082F]=8'hC1;
    mem['h0830]=8'hE5; mem['h0831]=8'hCD; mem['h0832]=8'h77; mem['h0833]=8'h0A;
    mem['h0834]=8'h22; mem['h0835]=8'h0C; mem['h0836]=8'h81; mem['h0837]=8'h21;
    mem['h0838]=8'h02; mem['h0839]=8'h00; mem['h083A]=8'h39; mem['h083B]=8'hCD;
    mem['h083C]=8'h35; mem['h083D]=8'h04; mem['h083E]=8'hD1; mem['h083F]=8'hC2;
    mem['h0840]=8'h57; mem['h0841]=8'h08; mem['h0842]=8'h09; mem['h0843]=8'hD5;
    mem['h0844]=8'h2B; mem['h0845]=8'h56; mem['h0846]=8'h2B; mem['h0847]=8'h5E;
    mem['h0848]=8'h23; mem['h0849]=8'h23; mem['h084A]=8'hE5; mem['h084B]=8'h2A;
    mem['h084C]=8'h0C; mem['h084D]=8'h81; mem['h084E]=8'hCD; mem['h084F]=8'h50;
    mem['h0850]=8'h07; mem['h0851]=8'hE1; mem['h0852]=8'hC2; mem['h0853]=8'h3B;
    mem['h0854]=8'h08; mem['h0855]=8'hD1; mem['h0856]=8'hF9; mem['h0857]=8'hEB;
    mem['h0858]=8'h0E; mem['h0859]=8'h08; mem['h085A]=8'hCD; mem['h085B]=8'h65;
    mem['h085C]=8'h04; mem['h085D]=8'hE5; mem['h085E]=8'h2A; mem['h085F]=8'h0C;
    mem['h0860]=8'h81; mem['h0861]=8'hE3; mem['h0862]=8'hE5; mem['h0863]=8'h2A;
    mem['h0864]=8'hA1; mem['h0865]=8'h80; mem['h0866]=8'hE3; mem['h0867]=8'hCD;
    mem['h0868]=8'h50; mem['h0869]=8'h0D; mem['h086A]=8'hCD; mem['h086B]=8'h56;
    mem['h086C]=8'h07; mem['h086D]=8'hA6; mem['h086E]=8'hCD; mem['h086F]=8'h4D;
    mem['h0870]=8'h0D; mem['h0871]=8'hE5; mem['h0872]=8'hCD; mem['h0873]=8'h7B;
    mem['h0874]=8'h17; mem['h0875]=8'hE1; mem['h0876]=8'hC5; mem['h0877]=8'hD5;
    mem['h0878]=8'h01; mem['h0879]=8'h00; mem['h087A]=8'h81; mem['h087B]=8'h51;
    mem['h087C]=8'h5A; mem['h087D]=8'h7E; mem['h087E]=8'hFE; mem['h087F]=8'hAB;
    mem['h0880]=8'h3E; mem['h0881]=8'h01; mem['h0882]=8'hC2; mem['h0883]=8'h93;
    mem['h0884]=8'h08; mem['h0885]=8'hCD; mem['h0886]=8'hE0; mem['h0887]=8'h08;
    mem['h0888]=8'hCD; mem['h0889]=8'h4D; mem['h088A]=8'h0D; mem['h088B]=8'hE5;
    mem['h088C]=8'hCD; mem['h088D]=8'h7B; mem['h088E]=8'h17; mem['h088F]=8'hCD;
    mem['h0890]=8'h2F; mem['h0891]=8'h17; mem['h0892]=8'hE1; mem['h0893]=8'hC5;
    mem['h0894]=8'hD5; mem['h0895]=8'hF5; mem['h0896]=8'h33; mem['h0897]=8'hE5;
    mem['h0898]=8'h2A; mem['h0899]=8'h13; mem['h089A]=8'h81; mem['h089B]=8'hE3;
    mem['h089C]=8'h06; mem['h089D]=8'h81; mem['h089E]=8'hC5; mem['h089F]=8'h33;
    mem['h08A0]=8'hCD; mem['h08A1]=8'h0B; mem['h08A2]=8'h09; mem['h08A3]=8'h22;
    mem['h08A4]=8'h13; mem['h08A5]=8'h81; mem['h08A6]=8'h7E; mem['h08A7]=8'hFE;
    mem['h08A8]=8'h3A; mem['h08A9]=8'hCA; mem['h08AA]=8'hC0; mem['h08AB]=8'h08;
    mem['h08AC]=8'hB7; mem['h08AD]=8'hC2; mem['h08AE]=8'h88; mem['h08AF]=8'h04;
    mem['h08B0]=8'h23; mem['h08B1]=8'h7E; mem['h08B2]=8'h23; mem['h08B3]=8'hB6;
    mem['h08B4]=8'hCA; mem['h08B5]=8'h32; mem['h08B6]=8'h09; mem['h08B7]=8'h23;
    mem['h08B8]=8'h5E; mem['h08B9]=8'h23; mem['h08BA]=8'h56; mem['h08BB]=8'hEB;
    mem['h08BC]=8'h22; mem['h08BD]=8'hA1; mem['h08BE]=8'h80; mem['h08BF]=8'hEB;
    mem['h08C0]=8'hCD; mem['h08C1]=8'hE0; mem['h08C2]=8'h08; mem['h08C3]=8'h11;
    mem['h08C4]=8'hA0; mem['h08C5]=8'h08; mem['h08C6]=8'hD5; mem['h08C7]=8'hC8;
    mem['h08C8]=8'hD6; mem['h08C9]=8'h80; mem['h08CA]=8'hDA; mem['h08CB]=8'h8E;
    mem['h08CC]=8'h0A; mem['h08CD]=8'hFE; mem['h08CE]=8'h25; mem['h08CF]=8'hD2;
    mem['h08D0]=8'h88; mem['h08D1]=8'h04; mem['h08D2]=8'h07; mem['h08D3]=8'h4F;
    mem['h08D4]=8'h06; mem['h08D5]=8'h00; mem['h08D6]=8'hEB; mem['h08D7]=8'h21;
    mem['h08D8]=8'h30; mem['h08D9]=8'h03; mem['h08DA]=8'h09; mem['h08DB]=8'h4E;
    mem['h08DC]=8'h23; mem['h08DD]=8'h46; mem['h08DE]=8'hC5; mem['h08DF]=8'hEB;
    mem['h08E0]=8'h23; mem['h08E1]=8'h7E; mem['h08E2]=8'hFE; mem['h08E3]=8'h3A;
    mem['h08E4]=8'hD0; mem['h08E5]=8'hFE; mem['h08E6]=8'h20; mem['h08E7]=8'hCA;
    mem['h08E8]=8'hE0; mem['h08E9]=8'h08; mem['h08EA]=8'hFE; mem['h08EB]=8'h30;
    mem['h08EC]=8'h3F; mem['h08ED]=8'h3C; mem['h08EE]=8'h3D; mem['h08EF]=8'hC9;
    mem['h08F0]=8'hEB; mem['h08F1]=8'h2A; mem['h08F2]=8'hA3; mem['h08F3]=8'h80;
    mem['h08F4]=8'hCA; mem['h08F5]=8'h05; mem['h08F6]=8'h09; mem['h08F7]=8'hEB;
    mem['h08F8]=8'hCD; mem['h08F9]=8'hAC; mem['h08FA]=8'h09; mem['h08FB]=8'hE5;
    mem['h08FC]=8'hCD; mem['h08FD]=8'h74; mem['h08FE]=8'h05; mem['h08FF]=8'h60;
    mem['h0900]=8'h69; mem['h0901]=8'hD1; mem['h0902]=8'hD2; mem['h0903]=8'h4D;
    mem['h0904]=8'h0A; mem['h0905]=8'h2B; mem['h0906]=8'h22; mem['h0907]=8'h21;
    mem['h0908]=8'h81; mem['h0909]=8'hEB; mem['h090A]=8'hC9; mem['h090B]=8'hDF;
    mem['h090C]=8'hC8; mem['h090D]=8'hD7; mem['h090E]=8'hFE; mem['h090F]=8'h1B;
    mem['h0910]=8'h28; mem['h0911]=8'h11; mem['h0912]=8'hFE; mem['h0913]=8'h03;
    mem['h0914]=8'h28; mem['h0915]=8'h0D; mem['h0916]=8'hFE; mem['h0917]=8'h13;
    mem['h0918]=8'hC0; mem['h0919]=8'hD7; mem['h091A]=8'hFE; mem['h091B]=8'h11;
    mem['h091C]=8'hC8; mem['h091D]=8'hFE; mem['h091E]=8'h03; mem['h091F]=8'h28;
    mem['h0920]=8'h07; mem['h0921]=8'h18; mem['h0922]=8'hF6; mem['h0923]=8'h3E;
    mem['h0924]=8'hFF; mem['h0925]=8'h32; mem['h0926]=8'h92; mem['h0927]=8'h80;
    mem['h0928]=8'hC0; mem['h0929]=8'hF6; mem['h092A]=8'hC0; mem['h092B]=8'h22;
    mem['h092C]=8'h13; mem['h092D]=8'h81; mem['h092E]=8'h21; mem['h092F]=8'hF6;
    mem['h0930]=8'hFF; mem['h0931]=8'hC1; mem['h0932]=8'h2A; mem['h0933]=8'hA1;
    mem['h0934]=8'h80; mem['h0935]=8'hF5; mem['h0936]=8'h7D; mem['h0937]=8'hA4;
    mem['h0938]=8'h3C; mem['h0939]=8'hCA; mem['h093A]=8'h45; mem['h093B]=8'h09;
    mem['h093C]=8'h22; mem['h093D]=8'h17; mem['h093E]=8'h81; mem['h093F]=8'h2A;
    mem['h0940]=8'h13; mem['h0941]=8'h81; mem['h0942]=8'h22; mem['h0943]=8'h19;
    mem['h0944]=8'h81; mem['h0945]=8'hAF; mem['h0946]=8'h32; mem['h0947]=8'h8A;
    mem['h0948]=8'h80; mem['h0949]=8'hCD; mem['h094A]=8'h7B; mem['h094B]=8'h0B;
    mem['h094C]=8'hF1; mem['h094D]=8'h21; mem['h094E]=8'h2B; mem['h094F]=8'h04;
    mem['h0950]=8'hC2; mem['h0951]=8'hBC; mem['h0952]=8'h04; mem['h0953]=8'hC3;
    mem['h0954]=8'hD3; mem['h0955]=8'h04; mem['h0956]=8'h2A; mem['h0957]=8'h19;
    mem['h0958]=8'h81; mem['h0959]=8'h7C; mem['h095A]=8'hB5; mem['h095B]=8'h1E;
    mem['h095C]=8'h20; mem['h095D]=8'hCA; mem['h095E]=8'h9C; mem['h095F]=8'h04;
    mem['h0960]=8'hEB; mem['h0961]=8'h2A; mem['h0962]=8'h17; mem['h0963]=8'h81;
    mem['h0964]=8'h22; mem['h0965]=8'hA1; mem['h0966]=8'h80; mem['h0967]=8'hEB;
    mem['h0968]=8'hC9; mem['h0969]=8'hCD; mem['h096A]=8'hAE; mem['h096B]=8'h14;
    mem['h096C]=8'hC0; mem['h096D]=8'h32; mem['h096E]=8'h86; mem['h096F]=8'h80;
    mem['h0970]=8'hC9; mem['h0971]=8'hE5; mem['h0972]=8'h2A; mem['h0973]=8'h8F;
    mem['h0974]=8'h80; mem['h0975]=8'h06; mem['h0976]=8'h00; mem['h0977]=8'h4F;
    mem['h0978]=8'h09; mem['h0979]=8'h22; mem['h097A]=8'h8F; mem['h097B]=8'h80;
    mem['h097C]=8'hE1; mem['h097D]=8'hC9; mem['h097E]=8'h7E; mem['h097F]=8'hFE;
    mem['h0980]=8'h41; mem['h0981]=8'hD8; mem['h0982]=8'hFE; mem['h0983]=8'h5B;
    mem['h0984]=8'h3F; mem['h0985]=8'hC9; mem['h0986]=8'hCD; mem['h0987]=8'hE0;
    mem['h0988]=8'h08; mem['h0989]=8'hCD; mem['h098A]=8'h4D; mem['h098B]=8'h0D;
    mem['h098C]=8'hCD; mem['h098D]=8'h2F; mem['h098E]=8'h17; mem['h098F]=8'hFA;
    mem['h0990]=8'hA7; mem['h0991]=8'h09; mem['h0992]=8'h3A; mem['h0993]=8'h2C;
    mem['h0994]=8'h81; mem['h0995]=8'hFE; mem['h0996]=8'h90; mem['h0997]=8'hDA;
    mem['h0998]=8'hD7; mem['h0999]=8'h17; mem['h099A]=8'h01; mem['h099B]=8'h80;
    mem['h099C]=8'h90; mem['h099D]=8'h11; mem['h099E]=8'h00; mem['h099F]=8'h00;
    mem['h09A0]=8'hE5; mem['h09A1]=8'hCD; mem['h09A2]=8'hAA; mem['h09A3]=8'h17;
    mem['h09A4]=8'hE1; mem['h09A5]=8'h51; mem['h09A6]=8'hC8; mem['h09A7]=8'h1E;
    mem['h09A8]=8'h08; mem['h09A9]=8'hC3; mem['h09AA]=8'h9C; mem['h09AB]=8'h04;
    mem['h09AC]=8'h2B; mem['h09AD]=8'h11; mem['h09AE]=8'h00; mem['h09AF]=8'h00;
    mem['h09B0]=8'hCD; mem['h09B1]=8'hE0; mem['h09B2]=8'h08; mem['h09B3]=8'hD0;
    mem['h09B4]=8'hE5; mem['h09B5]=8'hF5; mem['h09B6]=8'h21; mem['h09B7]=8'h98;
    mem['h09B8]=8'h19; mem['h09B9]=8'hCD; mem['h09BA]=8'h50; mem['h09BB]=8'h07;
    mem['h09BC]=8'hDA; mem['h09BD]=8'h88; mem['h09BE]=8'h04; mem['h09BF]=8'h62;
    mem['h09C0]=8'h6B; mem['h09C1]=8'h19; mem['h09C2]=8'h29; mem['h09C3]=8'h19;
    mem['h09C4]=8'h29; mem['h09C5]=8'hF1; mem['h09C6]=8'hD6; mem['h09C7]=8'h30;
    mem['h09C8]=8'h5F; mem['h09C9]=8'h16; mem['h09CA]=8'h00; mem['h09CB]=8'h19;
    mem['h09CC]=8'hEB; mem['h09CD]=8'hE1; mem['h09CE]=8'hC3; mem['h09CF]=8'hB0;
    mem['h09D0]=8'h09; mem['h09D1]=8'hCA; mem['h09D2]=8'hA4; mem['h09D3]=8'h05;
    mem['h09D4]=8'hCD; mem['h09D5]=8'h89; mem['h09D6]=8'h09; mem['h09D7]=8'h2B;
    mem['h09D8]=8'hCD; mem['h09D9]=8'hE0; mem['h09DA]=8'h08; mem['h09DB]=8'hE5;
    mem['h09DC]=8'h2A; mem['h09DD]=8'hF4; mem['h09DE]=8'h80; mem['h09DF]=8'hCA;
    mem['h09E0]=8'hF4; mem['h09E1]=8'h09; mem['h09E2]=8'hE1; mem['h09E3]=8'hCD;
    mem['h09E4]=8'h56; mem['h09E5]=8'h07; mem['h09E6]=8'h2C; mem['h09E7]=8'hD5;
    mem['h09E8]=8'hCD; mem['h09E9]=8'h89; mem['h09EA]=8'h09; mem['h09EB]=8'h2B;
    mem['h09EC]=8'hCD; mem['h09ED]=8'hE0; mem['h09EE]=8'h08; mem['h09EF]=8'hC2;
    mem['h09F0]=8'h88; mem['h09F1]=8'h04; mem['h09F2]=8'hE3; mem['h09F3]=8'hEB;
    mem['h09F4]=8'h7D; mem['h09F5]=8'h93; mem['h09F6]=8'h5F; mem['h09F7]=8'h7C;
    mem['h09F8]=8'h9A; mem['h09F9]=8'h57; mem['h09FA]=8'hDA; mem['h09FB]=8'h7D;
    mem['h09FC]=8'h04; mem['h09FD]=8'hE5; mem['h09FE]=8'h2A; mem['h09FF]=8'h1B;
    mem['h0A00]=8'h81; mem['h0A01]=8'h01; mem['h0A02]=8'h28; mem['h0A03]=8'h00;
    mem['h0A04]=8'h09; mem['h0A05]=8'hCD; mem['h0A06]=8'h50; mem['h0A07]=8'h07;
    mem['h0A08]=8'hD2; mem['h0A09]=8'h7D; mem['h0A0A]=8'h04; mem['h0A0B]=8'hEB;
    mem['h0A0C]=8'h22; mem['h0A0D]=8'h9F; mem['h0A0E]=8'h80; mem['h0A0F]=8'hE1;
    mem['h0A10]=8'h22; mem['h0A11]=8'hF4; mem['h0A12]=8'h80; mem['h0A13]=8'hE1;
    mem['h0A14]=8'hC3; mem['h0A15]=8'hA4; mem['h0A16]=8'h05; mem['h0A17]=8'hCA;
    mem['h0A18]=8'hA0; mem['h0A19]=8'h05; mem['h0A1A]=8'hCD; mem['h0A1B]=8'hA4;
    mem['h0A1C]=8'h05; mem['h0A1D]=8'h01; mem['h0A1E]=8'hA0; mem['h0A1F]=8'h08;
    mem['h0A20]=8'hC3; mem['h0A21]=8'h33; mem['h0A22]=8'h0A; mem['h0A23]=8'h0E;
    mem['h0A24]=8'h03; mem['h0A25]=8'hCD; mem['h0A26]=8'h65; mem['h0A27]=8'h04;
    mem['h0A28]=8'hC1; mem['h0A29]=8'hE5; mem['h0A2A]=8'hE5; mem['h0A2B]=8'h2A;
    mem['h0A2C]=8'hA1; mem['h0A2D]=8'h80; mem['h0A2E]=8'hE3; mem['h0A2F]=8'h3E;
    mem['h0A30]=8'h8C; mem['h0A31]=8'hF5; mem['h0A32]=8'h33; mem['h0A33]=8'hC5;
    mem['h0A34]=8'hCD; mem['h0A35]=8'hAC; mem['h0A36]=8'h09; mem['h0A37]=8'hCD;
    mem['h0A38]=8'h79; mem['h0A39]=8'h0A; mem['h0A3A]=8'hE5; mem['h0A3B]=8'h2A;
    mem['h0A3C]=8'hA1; mem['h0A3D]=8'h80; mem['h0A3E]=8'hCD; mem['h0A3F]=8'h50;
    mem['h0A40]=8'h07; mem['h0A41]=8'hE1; mem['h0A42]=8'h23; mem['h0A43]=8'hDC;
    mem['h0A44]=8'h77; mem['h0A45]=8'h05; mem['h0A46]=8'hD4; mem['h0A47]=8'h74;
    mem['h0A48]=8'h05; mem['h0A49]=8'h60; mem['h0A4A]=8'h69; mem['h0A4B]=8'h2B;
    mem['h0A4C]=8'hD8; mem['h0A4D]=8'h1E; mem['h0A4E]=8'h0E; mem['h0A4F]=8'hC3;
    mem['h0A50]=8'h9C; mem['h0A51]=8'h04; mem['h0A52]=8'hC0; mem['h0A53]=8'h16;
    mem['h0A54]=8'hFF; mem['h0A55]=8'hCD; mem['h0A56]=8'h31; mem['h0A57]=8'h04;
    mem['h0A58]=8'hF9; mem['h0A59]=8'hFE; mem['h0A5A]=8'h8C; mem['h0A5B]=8'h1E;
    mem['h0A5C]=8'h04; mem['h0A5D]=8'hC2; mem['h0A5E]=8'h9C; mem['h0A5F]=8'h04;
    mem['h0A60]=8'hE1; mem['h0A61]=8'h22; mem['h0A62]=8'hA1; mem['h0A63]=8'h80;
    mem['h0A64]=8'h23; mem['h0A65]=8'h7C; mem['h0A66]=8'hB5; mem['h0A67]=8'hC2;
    mem['h0A68]=8'h71; mem['h0A69]=8'h0A; mem['h0A6A]=8'h3A; mem['h0A6B]=8'h11;
    mem['h0A6C]=8'h81; mem['h0A6D]=8'hB7; mem['h0A6E]=8'hC2; mem['h0A6F]=8'hD2;
    mem['h0A70]=8'h04; mem['h0A71]=8'h21; mem['h0A72]=8'hA0; mem['h0A73]=8'h08;
    mem['h0A74]=8'hE3; mem['h0A75]=8'h3E; mem['h0A76]=8'hE1; mem['h0A77]=8'h01;
    mem['h0A78]=8'h3A; mem['h0A79]=8'h0E; mem['h0A7A]=8'h00; mem['h0A7B]=8'h06;
    mem['h0A7C]=8'h00; mem['h0A7D]=8'h79; mem['h0A7E]=8'h48; mem['h0A7F]=8'h47;
    mem['h0A80]=8'h7E; mem['h0A81]=8'hB7; mem['h0A82]=8'hC8; mem['h0A83]=8'hB8;
    mem['h0A84]=8'hC8; mem['h0A85]=8'h23; mem['h0A86]=8'hFE; mem['h0A87]=8'h22;
    mem['h0A88]=8'hCA; mem['h0A89]=8'h7D; mem['h0A8A]=8'h0A; mem['h0A8B]=8'hC3;
    mem['h0A8C]=8'h80; mem['h0A8D]=8'h0A; mem['h0A8E]=8'hCD; mem['h0A8F]=8'h43;
    mem['h0A90]=8'h0F; mem['h0A91]=8'hCD; mem['h0A92]=8'h56; mem['h0A93]=8'h07;
    mem['h0A94]=8'hB4; mem['h0A95]=8'hD5; mem['h0A96]=8'h3A; mem['h0A97]=8'hF2;
    mem['h0A98]=8'h80; mem['h0A99]=8'hF5; mem['h0A9A]=8'hCD; mem['h0A9B]=8'h5F;
    mem['h0A9C]=8'h0D; mem['h0A9D]=8'hF1; mem['h0A9E]=8'hE3; mem['h0A9F]=8'h22;
    mem['h0AA0]=8'h13; mem['h0AA1]=8'h81; mem['h0AA2]=8'h1F; mem['h0AA3]=8'hCD;
    mem['h0AA4]=8'h52; mem['h0AA5]=8'h0D; mem['h0AA6]=8'hCA; mem['h0AA7]=8'hE1;
    mem['h0AA8]=8'h0A; mem['h0AA9]=8'hE5; mem['h0AAA]=8'h2A; mem['h0AAB]=8'h29;
    mem['h0AAC]=8'h81; mem['h0AAD]=8'hE5; mem['h0AAE]=8'h23; mem['h0AAF]=8'h23;
    mem['h0AB0]=8'h5E; mem['h0AB1]=8'h23; mem['h0AB2]=8'h56; mem['h0AB3]=8'h2A;
    mem['h0AB4]=8'hA3; mem['h0AB5]=8'h80; mem['h0AB6]=8'hCD; mem['h0AB7]=8'h50;
    mem['h0AB8]=8'h07; mem['h0AB9]=8'hD2; mem['h0ABA]=8'hD0; mem['h0ABB]=8'h0A;
    mem['h0ABC]=8'h2A; mem['h0ABD]=8'h9F; mem['h0ABE]=8'h80; mem['h0ABF]=8'hCD;
    mem['h0AC0]=8'h50; mem['h0AC1]=8'h07; mem['h0AC2]=8'hD1; mem['h0AC3]=8'hD2;
    mem['h0AC4]=8'hD8; mem['h0AC5]=8'h0A; mem['h0AC6]=8'h21; mem['h0AC7]=8'h04;
    mem['h0AC8]=8'h81; mem['h0AC9]=8'hCD; mem['h0ACA]=8'h50; mem['h0ACB]=8'h07;
    mem['h0ACC]=8'hD2; mem['h0ACD]=8'hD8; mem['h0ACE]=8'h0A; mem['h0ACF]=8'h3E;
    mem['h0AD0]=8'hD1; mem['h0AD1]=8'hCD; mem['h0AD2]=8'h87; mem['h0AD3]=8'h13;
    mem['h0AD4]=8'hEB; mem['h0AD5]=8'hCD; mem['h0AD6]=8'hC0; mem['h0AD7]=8'h11;
    mem['h0AD8]=8'hCD; mem['h0AD9]=8'h87; mem['h0ADA]=8'h13; mem['h0ADB]=8'hE1;
    mem['h0ADC]=8'hCD; mem['h0ADD]=8'h8A; mem['h0ADE]=8'h17; mem['h0ADF]=8'hE1;
    mem['h0AE0]=8'hC9; mem['h0AE1]=8'hE5; mem['h0AE2]=8'hCD; mem['h0AE3]=8'h87;
    mem['h0AE4]=8'h17; mem['h0AE5]=8'hD1; mem['h0AE6]=8'hE1; mem['h0AE7]=8'hC9;
    mem['h0AE8]=8'hCD; mem['h0AE9]=8'hAE; mem['h0AEA]=8'h14; mem['h0AEB]=8'h7E;
    mem['h0AEC]=8'h47; mem['h0AED]=8'hFE; mem['h0AEE]=8'h8C; mem['h0AEF]=8'hCA;
    mem['h0AF0]=8'hF7; mem['h0AF1]=8'h0A; mem['h0AF2]=8'hCD; mem['h0AF3]=8'h56;
    mem['h0AF4]=8'h07; mem['h0AF5]=8'h88; mem['h0AF6]=8'h2B; mem['h0AF7]=8'h4B;
    mem['h0AF8]=8'h0D; mem['h0AF9]=8'h78; mem['h0AFA]=8'hCA; mem['h0AFB]=8'hC8;
    mem['h0AFC]=8'h08; mem['h0AFD]=8'hCD; mem['h0AFE]=8'hAD; mem['h0AFF]=8'h09;
    mem['h0B00]=8'hFE; mem['h0B01]=8'h2C; mem['h0B02]=8'hC0; mem['h0B03]=8'hC3;
    mem['h0B04]=8'hF8; mem['h0B05]=8'h0A; mem['h0B06]=8'hCD; mem['h0B07]=8'h5F;
    mem['h0B08]=8'h0D; mem['h0B09]=8'h7E; mem['h0B0A]=8'hFE; mem['h0B0B]=8'h88;
    mem['h0B0C]=8'hCA; mem['h0B0D]=8'h14; mem['h0B0E]=8'h0B; mem['h0B0F]=8'hCD;
    mem['h0B10]=8'h56; mem['h0B11]=8'h07; mem['h0B12]=8'hA9; mem['h0B13]=8'h2B;
    mem['h0B14]=8'hCD; mem['h0B15]=8'h50; mem['h0B16]=8'h0D; mem['h0B17]=8'hCD;
    mem['h0B18]=8'h2F; mem['h0B19]=8'h17; mem['h0B1A]=8'hCA; mem['h0B1B]=8'h79;
    mem['h0B1C]=8'h0A; mem['h0B1D]=8'hCD; mem['h0B1E]=8'hE0; mem['h0B1F]=8'h08;
    mem['h0B20]=8'hDA; mem['h0B21]=8'h34; mem['h0B22]=8'h0A; mem['h0B23]=8'hC3;
    mem['h0B24]=8'hC7; mem['h0B25]=8'h08; mem['h0B26]=8'h2B; mem['h0B27]=8'hCD;
    mem['h0B28]=8'hE0; mem['h0B29]=8'h08; mem['h0B2A]=8'hCA; mem['h0B2B]=8'h88;
    mem['h0B2C]=8'h0B; mem['h0B2D]=8'hC8; mem['h0B2E]=8'hFE; mem['h0B2F]=8'hA5;
    mem['h0B30]=8'hCA; mem['h0B31]=8'hBB; mem['h0B32]=8'h0B; mem['h0B33]=8'hFE;
    mem['h0B34]=8'hA8; mem['h0B35]=8'hCA; mem['h0B36]=8'hBB; mem['h0B37]=8'h0B;
    mem['h0B38]=8'hE5; mem['h0B39]=8'hFE; mem['h0B3A]=8'h2C; mem['h0B3B]=8'hCA;
    mem['h0B3C]=8'hA4; mem['h0B3D]=8'h0B; mem['h0B3E]=8'hFE; mem['h0B3F]=8'h3B;
    mem['h0B40]=8'hCA; mem['h0B41]=8'hDE; mem['h0B42]=8'h0B; mem['h0B43]=8'hC1;
    mem['h0B44]=8'hCD; mem['h0B45]=8'h5F; mem['h0B46]=8'h0D; mem['h0B47]=8'hE5;
    mem['h0B48]=8'h3A; mem['h0B49]=8'hF2; mem['h0B4A]=8'h80; mem['h0B4B]=8'hB7;
    mem['h0B4C]=8'hC2; mem['h0B4D]=8'h74; mem['h0B4E]=8'h0B; mem['h0B4F]=8'hCD;
    mem['h0B50]=8'hD4; mem['h0B51]=8'h18; mem['h0B52]=8'hCD; mem['h0B53]=8'hE4;
    mem['h0B54]=8'h11; mem['h0B55]=8'h36; mem['h0B56]=8'h20; mem['h0B57]=8'h2A;
    mem['h0B58]=8'h29; mem['h0B59]=8'h81; mem['h0B5A]=8'h34; mem['h0B5B]=8'h2A;
    mem['h0B5C]=8'h29; mem['h0B5D]=8'h81; mem['h0B5E]=8'h3A; mem['h0B5F]=8'h87;
    mem['h0B60]=8'h80; mem['h0B61]=8'h47; mem['h0B62]=8'h04; mem['h0B63]=8'hCA;
    mem['h0B64]=8'h70; mem['h0B65]=8'h0B; mem['h0B66]=8'h04; mem['h0B67]=8'h3A;
    mem['h0B68]=8'hF0; mem['h0B69]=8'h80; mem['h0B6A]=8'h86; mem['h0B6B]=8'h3D;
    mem['h0B6C]=8'hB8; mem['h0B6D]=8'hD4; mem['h0B6E]=8'h88; mem['h0B6F]=8'h0B;
    mem['h0B70]=8'hCD; mem['h0B71]=8'h29; mem['h0B72]=8'h12; mem['h0B73]=8'hAF;
    mem['h0B74]=8'hC4; mem['h0B75]=8'h29; mem['h0B76]=8'h12; mem['h0B77]=8'hE1;
    mem['h0B78]=8'hC3; mem['h0B79]=8'h26; mem['h0B7A]=8'h0B; mem['h0B7B]=8'h3A;
    mem['h0B7C]=8'hF0; mem['h0B7D]=8'h80; mem['h0B7E]=8'hB7; mem['h0B7F]=8'hC8;
    mem['h0B80]=8'hC3; mem['h0B81]=8'h88; mem['h0B82]=8'h0B; mem['h0B83]=8'h36;
    mem['h0B84]=8'h00; mem['h0B85]=8'h21; mem['h0B86]=8'hA5; mem['h0B87]=8'h80;
    mem['h0B88]=8'h3E; mem['h0B89]=8'h0D; mem['h0B8A]=8'hCD; mem['h0B8B]=8'h61;
    mem['h0B8C]=8'h07; mem['h0B8D]=8'h3E; mem['h0B8E]=8'h0A; mem['h0B8F]=8'hCD;
    mem['h0B90]=8'h61; mem['h0B91]=8'h07; mem['h0B92]=8'hAF; mem['h0B93]=8'h32;
    mem['h0B94]=8'hF0; mem['h0B95]=8'h80; mem['h0B96]=8'h3A; mem['h0B97]=8'h86;
    mem['h0B98]=8'h80; mem['h0B99]=8'h3D; mem['h0B9A]=8'hC8; mem['h0B9B]=8'hF5;
    mem['h0B9C]=8'hAF; mem['h0B9D]=8'hCD; mem['h0B9E]=8'h61; mem['h0B9F]=8'h07;
    mem['h0BA0]=8'hF1; mem['h0BA1]=8'hC3; mem['h0BA2]=8'h99; mem['h0BA3]=8'h0B;
    mem['h0BA4]=8'h3A; mem['h0BA5]=8'h88; mem['h0BA6]=8'h80; mem['h0BA7]=8'h47;
    mem['h0BA8]=8'h3A; mem['h0BA9]=8'hF0; mem['h0BAA]=8'h80; mem['h0BAB]=8'hB8;
    mem['h0BAC]=8'hD4; mem['h0BAD]=8'h88; mem['h0BAE]=8'h0B; mem['h0BAF]=8'hD2;
    mem['h0BB0]=8'hDE; mem['h0BB1]=8'h0B; mem['h0BB2]=8'hD6; mem['h0BB3]=8'h0E;
    mem['h0BB4]=8'hD2; mem['h0BB5]=8'hB2; mem['h0BB6]=8'h0B; mem['h0BB7]=8'h2F;
    mem['h0BB8]=8'hC3; mem['h0BB9]=8'hD3; mem['h0BBA]=8'h0B; mem['h0BBB]=8'hF5;
    mem['h0BBC]=8'hCD; mem['h0BBD]=8'hAB; mem['h0BBE]=8'h14; mem['h0BBF]=8'hCD;
    mem['h0BC0]=8'h56; mem['h0BC1]=8'h07; mem['h0BC2]=8'h29; mem['h0BC3]=8'h2B;
    mem['h0BC4]=8'hF1; mem['h0BC5]=8'hD6; mem['h0BC6]=8'hA8; mem['h0BC7]=8'hE5;
    mem['h0BC8]=8'hCA; mem['h0BC9]=8'hCE; mem['h0BCA]=8'h0B; mem['h0BCB]=8'h3A;
    mem['h0BCC]=8'hF0; mem['h0BCD]=8'h80; mem['h0BCE]=8'h2F; mem['h0BCF]=8'h83;
    mem['h0BD0]=8'hD2; mem['h0BD1]=8'hDE; mem['h0BD2]=8'h0B; mem['h0BD3]=8'h3C;
    mem['h0BD4]=8'h47; mem['h0BD5]=8'h3E; mem['h0BD6]=8'h20; mem['h0BD7]=8'hCD;
    mem['h0BD8]=8'h61; mem['h0BD9]=8'h07; mem['h0BDA]=8'h05; mem['h0BDB]=8'hC2;
    mem['h0BDC]=8'hD7; mem['h0BDD]=8'h0B; mem['h0BDE]=8'hE1; mem['h0BDF]=8'hCD;
    mem['h0BE0]=8'hE0; mem['h0BE1]=8'h08; mem['h0BE2]=8'hC3; mem['h0BE3]=8'h2D;
    mem['h0BE4]=8'h0B; mem['h0BE5]=8'h3F; mem['h0BE6]=8'h52; mem['h0BE7]=8'h65;
    mem['h0BE8]=8'h64; mem['h0BE9]=8'h6F; mem['h0BEA]=8'h20; mem['h0BEB]=8'h66;
    mem['h0BEC]=8'h72; mem['h0BED]=8'h6F; mem['h0BEE]=8'h6D; mem['h0BEF]=8'h20;
    mem['h0BF0]=8'h73; mem['h0BF1]=8'h74; mem['h0BF2]=8'h61; mem['h0BF3]=8'h72;
    mem['h0BF4]=8'h74; mem['h0BF5]=8'h0D; mem['h0BF6]=8'h0A; mem['h0BF7]=8'h00;
    mem['h0BF8]=8'h3A; mem['h0BF9]=8'h12; mem['h0BFA]=8'h81; mem['h0BFB]=8'hB7;
    mem['h0BFC]=8'hC2; mem['h0BFD]=8'h82; mem['h0BFE]=8'h04; mem['h0BFF]=8'hC1;
    mem['h0C00]=8'h21; mem['h0C01]=8'hE5; mem['h0C02]=8'h0B; mem['h0C03]=8'hCD;
    mem['h0C04]=8'h26; mem['h0C05]=8'h12; mem['h0C06]=8'hC3; mem['h0C07]=8'hD3;
    mem['h0C08]=8'h05; mem['h0C09]=8'hCD; mem['h0C0A]=8'h91; mem['h0C0B]=8'h11;
    mem['h0C0C]=8'h7E; mem['h0C0D]=8'hFE; mem['h0C0E]=8'h22; mem['h0C0F]=8'h3E;
    mem['h0C10]=8'h00; mem['h0C11]=8'h32; mem['h0C12]=8'h8A; mem['h0C13]=8'h80;
    mem['h0C14]=8'hC2; mem['h0C15]=8'h23; mem['h0C16]=8'h0C; mem['h0C17]=8'hCD;
    mem['h0C18]=8'hE5; mem['h0C19]=8'h11; mem['h0C1A]=8'hCD; mem['h0C1B]=8'h56;
    mem['h0C1C]=8'h07; mem['h0C1D]=8'h3B; mem['h0C1E]=8'hE5; mem['h0C1F]=8'hCD;
    mem['h0C20]=8'h29; mem['h0C21]=8'h12; mem['h0C22]=8'h3E; mem['h0C23]=8'hE5;
    mem['h0C24]=8'hCD; mem['h0C25]=8'hD7; mem['h0C26]=8'h05; mem['h0C27]=8'hC1;
    mem['h0C28]=8'hDA; mem['h0C29]=8'h2F; mem['h0C2A]=8'h09; mem['h0C2B]=8'h23;
    mem['h0C2C]=8'h7E; mem['h0C2D]=8'hB7; mem['h0C2E]=8'h2B; mem['h0C2F]=8'hC5;
    mem['h0C30]=8'hCA; mem['h0C31]=8'h76; mem['h0C32]=8'h0A; mem['h0C33]=8'h36;
    mem['h0C34]=8'h2C; mem['h0C35]=8'hC3; mem['h0C36]=8'h3D; mem['h0C37]=8'h0C;
    mem['h0C38]=8'hE5; mem['h0C39]=8'h2A; mem['h0C3A]=8'h21; mem['h0C3B]=8'h81;
    mem['h0C3C]=8'hF6; mem['h0C3D]=8'hAF; mem['h0C3E]=8'h32; mem['h0C3F]=8'h12;
    mem['h0C40]=8'h81; mem['h0C41]=8'hE3; mem['h0C42]=8'hC3; mem['h0C43]=8'h49;
    mem['h0C44]=8'h0C; mem['h0C45]=8'hCD; mem['h0C46]=8'h56; mem['h0C47]=8'h07;
    mem['h0C48]=8'h2C; mem['h0C49]=8'hCD; mem['h0C4A]=8'h43; mem['h0C4B]=8'h0F;
    mem['h0C4C]=8'hE3; mem['h0C4D]=8'hD5; mem['h0C4E]=8'h7E; mem['h0C4F]=8'hFE;
    mem['h0C50]=8'h2C; mem['h0C51]=8'hCA; mem['h0C52]=8'h71; mem['h0C53]=8'h0C;
    mem['h0C54]=8'h3A; mem['h0C55]=8'h12; mem['h0C56]=8'h81; mem['h0C57]=8'hB7;
    mem['h0C58]=8'hC2; mem['h0C59]=8'hDE; mem['h0C5A]=8'h0C; mem['h0C5B]=8'h3E;
    mem['h0C5C]=8'h3F; mem['h0C5D]=8'hCD; mem['h0C5E]=8'h61; mem['h0C5F]=8'h07;
    mem['h0C60]=8'hCD; mem['h0C61]=8'hD7; mem['h0C62]=8'h05; mem['h0C63]=8'hD1;
    mem['h0C64]=8'hC1; mem['h0C65]=8'hDA; mem['h0C66]=8'h2F; mem['h0C67]=8'h09;
    mem['h0C68]=8'h23; mem['h0C69]=8'h7E; mem['h0C6A]=8'hB7; mem['h0C6B]=8'h2B;
    mem['h0C6C]=8'hC5; mem['h0C6D]=8'hCA; mem['h0C6E]=8'h76; mem['h0C6F]=8'h0A;
    mem['h0C70]=8'hD5; mem['h0C71]=8'h3A; mem['h0C72]=8'hF2; mem['h0C73]=8'h80;
    mem['h0C74]=8'hB7; mem['h0C75]=8'hCA; mem['h0C76]=8'h9B; mem['h0C77]=8'h0C;
    mem['h0C78]=8'hCD; mem['h0C79]=8'hE0; mem['h0C7A]=8'h08; mem['h0C7B]=8'h57;
    mem['h0C7C]=8'h47; mem['h0C7D]=8'hFE; mem['h0C7E]=8'h22; mem['h0C7F]=8'hCA;
    mem['h0C80]=8'h8F; mem['h0C81]=8'h0C; mem['h0C82]=8'h3A; mem['h0C83]=8'h12;
    mem['h0C84]=8'h81; mem['h0C85]=8'hB7; mem['h0C86]=8'h57; mem['h0C87]=8'hCA;
    mem['h0C88]=8'h8C; mem['h0C89]=8'h0C; mem['h0C8A]=8'h16; mem['h0C8B]=8'h3A;
    mem['h0C8C]=8'h06; mem['h0C8D]=8'h2C; mem['h0C8E]=8'h2B; mem['h0C8F]=8'hCD;
    mem['h0C90]=8'hE8; mem['h0C91]=8'h11; mem['h0C92]=8'hEB; mem['h0C93]=8'h21;
    mem['h0C94]=8'hA6; mem['h0C95]=8'h0C; mem['h0C96]=8'hE3; mem['h0C97]=8'hD5;
    mem['h0C98]=8'hC3; mem['h0C99]=8'hA9; mem['h0C9A]=8'h0A; mem['h0C9B]=8'hCD;
    mem['h0C9C]=8'hE0; mem['h0C9D]=8'h08; mem['h0C9E]=8'hCD; mem['h0C9F]=8'h36;
    mem['h0CA0]=8'h18; mem['h0CA1]=8'hE3; mem['h0CA2]=8'hCD; mem['h0CA3]=8'h87;
    mem['h0CA4]=8'h17; mem['h0CA5]=8'hE1; mem['h0CA6]=8'h2B; mem['h0CA7]=8'hCD;
    mem['h0CA8]=8'hE0; mem['h0CA9]=8'h08; mem['h0CAA]=8'hCA; mem['h0CAB]=8'hB2;
    mem['h0CAC]=8'h0C; mem['h0CAD]=8'hFE; mem['h0CAE]=8'h2C; mem['h0CAF]=8'hC2;
    mem['h0CB0]=8'hF8; mem['h0CB1]=8'h0B; mem['h0CB2]=8'hE3; mem['h0CB3]=8'h2B;
    mem['h0CB4]=8'hCD; mem['h0CB5]=8'hE0; mem['h0CB6]=8'h08; mem['h0CB7]=8'hC2;
    mem['h0CB8]=8'h45; mem['h0CB9]=8'h0C; mem['h0CBA]=8'hD1; mem['h0CBB]=8'h3A;
    mem['h0CBC]=8'h12; mem['h0CBD]=8'h81; mem['h0CBE]=8'hB7; mem['h0CBF]=8'hEB;
    mem['h0CC0]=8'hC2; mem['h0CC1]=8'h06; mem['h0CC2]=8'h09; mem['h0CC3]=8'hD5;
    mem['h0CC4]=8'hB6; mem['h0CC5]=8'h21; mem['h0CC6]=8'hCD; mem['h0CC7]=8'h0C;
    mem['h0CC8]=8'hC4; mem['h0CC9]=8'h26; mem['h0CCA]=8'h12; mem['h0CCB]=8'hE1;
    mem['h0CCC]=8'hC9; mem['h0CCD]=8'h3F; mem['h0CCE]=8'h45; mem['h0CCF]=8'h78;
    mem['h0CD0]=8'h74; mem['h0CD1]=8'h72; mem['h0CD2]=8'h61; mem['h0CD3]=8'h20;
    mem['h0CD4]=8'h69; mem['h0CD5]=8'h67; mem['h0CD6]=8'h6E; mem['h0CD7]=8'h6F;
    mem['h0CD8]=8'h72; mem['h0CD9]=8'h65; mem['h0CDA]=8'h64; mem['h0CDB]=8'h0D;
    mem['h0CDC]=8'h0A; mem['h0CDD]=8'h00; mem['h0CDE]=8'hCD; mem['h0CDF]=8'h77;
    mem['h0CE0]=8'h0A; mem['h0CE1]=8'hB7; mem['h0CE2]=8'hC2; mem['h0CE3]=8'hF7;
    mem['h0CE4]=8'h0C; mem['h0CE5]=8'h23; mem['h0CE6]=8'h7E; mem['h0CE7]=8'h23;
    mem['h0CE8]=8'hB6; mem['h0CE9]=8'h1E; mem['h0CEA]=8'h06; mem['h0CEB]=8'hCA;
    mem['h0CEC]=8'h9C; mem['h0CED]=8'h04; mem['h0CEE]=8'h23; mem['h0CEF]=8'h5E;
    mem['h0CF0]=8'h23; mem['h0CF1]=8'h56; mem['h0CF2]=8'hEB; mem['h0CF3]=8'h22;
    mem['h0CF4]=8'h0E; mem['h0CF5]=8'h81; mem['h0CF6]=8'hEB; mem['h0CF7]=8'hCD;
    mem['h0CF8]=8'hE0; mem['h0CF9]=8'h08; mem['h0CFA]=8'hFE; mem['h0CFB]=8'h83;
    mem['h0CFC]=8'hC2; mem['h0CFD]=8'hDE; mem['h0CFE]=8'h0C; mem['h0CFF]=8'hC3;
    mem['h0D00]=8'h71; mem['h0D01]=8'h0C; mem['h0D02]=8'h11; mem['h0D03]=8'h00;
    mem['h0D04]=8'h00; mem['h0D05]=8'hC4; mem['h0D06]=8'h43; mem['h0D07]=8'h0F;
    mem['h0D08]=8'h22; mem['h0D09]=8'h13; mem['h0D0A]=8'h81; mem['h0D0B]=8'hCD;
    mem['h0D0C]=8'h31; mem['h0D0D]=8'h04; mem['h0D0E]=8'hC2; mem['h0D0F]=8'h8E;
    mem['h0D10]=8'h04; mem['h0D11]=8'hF9; mem['h0D12]=8'hD5; mem['h0D13]=8'h7E;
    mem['h0D14]=8'h23; mem['h0D15]=8'hF5; mem['h0D16]=8'hD5; mem['h0D17]=8'hCD;
    mem['h0D18]=8'h6D; mem['h0D19]=8'h17; mem['h0D1A]=8'hE3; mem['h0D1B]=8'hE5;
    mem['h0D1C]=8'hCD; mem['h0D1D]=8'hDA; mem['h0D1E]=8'h14; mem['h0D1F]=8'hE1;
    mem['h0D20]=8'hCD; mem['h0D21]=8'h87; mem['h0D22]=8'h17; mem['h0D23]=8'hE1;
    mem['h0D24]=8'hCD; mem['h0D25]=8'h7E; mem['h0D26]=8'h17; mem['h0D27]=8'hE5;
    mem['h0D28]=8'hCD; mem['h0D29]=8'hAA; mem['h0D2A]=8'h17; mem['h0D2B]=8'hE1;
    mem['h0D2C]=8'hC1; mem['h0D2D]=8'h90; mem['h0D2E]=8'hCD; mem['h0D2F]=8'h7E;
    mem['h0D30]=8'h17; mem['h0D31]=8'hCA; mem['h0D32]=8'h3D; mem['h0D33]=8'h0D;
    mem['h0D34]=8'hEB; mem['h0D35]=8'h22; mem['h0D36]=8'hA1; mem['h0D37]=8'h80;
    mem['h0D38]=8'h69; mem['h0D39]=8'h60; mem['h0D3A]=8'hC3; mem['h0D3B]=8'h9C;
    mem['h0D3C]=8'h08; mem['h0D3D]=8'hF9; mem['h0D3E]=8'h2A; mem['h0D3F]=8'h13;
    mem['h0D40]=8'h81; mem['h0D41]=8'h7E; mem['h0D42]=8'hFE; mem['h0D43]=8'h2C;
    mem['h0D44]=8'hC2; mem['h0D45]=8'hA0; mem['h0D46]=8'h08; mem['h0D47]=8'hCD;
    mem['h0D48]=8'hE0; mem['h0D49]=8'h08; mem['h0D4A]=8'hCD; mem['h0D4B]=8'h05;
    mem['h0D4C]=8'h0D; mem['h0D4D]=8'hCD; mem['h0D4E]=8'h5F; mem['h0D4F]=8'h0D;
    mem['h0D50]=8'hF6; mem['h0D51]=8'h37; mem['h0D52]=8'h3A; mem['h0D53]=8'hF2;
    mem['h0D54]=8'h80; mem['h0D55]=8'h8F; mem['h0D56]=8'hB7; mem['h0D57]=8'hE8;
    mem['h0D58]=8'hC3; mem['h0D59]=8'h9A; mem['h0D5A]=8'h04; mem['h0D5B]=8'hCD;
    mem['h0D5C]=8'h56; mem['h0D5D]=8'h07; mem['h0D5E]=8'h28; mem['h0D5F]=8'h2B;
    mem['h0D60]=8'h16; mem['h0D61]=8'h00; mem['h0D62]=8'hD5; mem['h0D63]=8'h0E;
    mem['h0D64]=8'h01; mem['h0D65]=8'hCD; mem['h0D66]=8'h65; mem['h0D67]=8'h04;
    mem['h0D68]=8'hCD; mem['h0D69]=8'hD6; mem['h0D6A]=8'h0D; mem['h0D6B]=8'h22;
    mem['h0D6C]=8'h15; mem['h0D6D]=8'h81; mem['h0D6E]=8'h2A; mem['h0D6F]=8'h15;
    mem['h0D70]=8'h81; mem['h0D71]=8'hC1; mem['h0D72]=8'h78; mem['h0D73]=8'hFE;
    mem['h0D74]=8'h78; mem['h0D75]=8'hD4; mem['h0D76]=8'h50; mem['h0D77]=8'h0D;
    mem['h0D78]=8'h7E; mem['h0D79]=8'h16; mem['h0D7A]=8'h00; mem['h0D7B]=8'hD6;
    mem['h0D7C]=8'hB3; mem['h0D7D]=8'hDA; mem['h0D7E]=8'h97; mem['h0D7F]=8'h0D;
    mem['h0D80]=8'hFE; mem['h0D81]=8'h03; mem['h0D82]=8'hD2; mem['h0D83]=8'h97;
    mem['h0D84]=8'h0D; mem['h0D85]=8'hFE; mem['h0D86]=8'h01; mem['h0D87]=8'h17;
    mem['h0D88]=8'hAA; mem['h0D89]=8'hBA; mem['h0D8A]=8'h57; mem['h0D8B]=8'hDA;
    mem['h0D8C]=8'h88; mem['h0D8D]=8'h04; mem['h0D8E]=8'h22; mem['h0D8F]=8'h0A;
    mem['h0D90]=8'h81; mem['h0D91]=8'hCD; mem['h0D92]=8'hE0; mem['h0D93]=8'h08;
    mem['h0D94]=8'hC3; mem['h0D95]=8'h7B; mem['h0D96]=8'h0D; mem['h0D97]=8'h7A;
    mem['h0D98]=8'hB7; mem['h0D99]=8'hC2; mem['h0D9A]=8'hBE; mem['h0D9B]=8'h0E;
    mem['h0D9C]=8'h7E; mem['h0D9D]=8'h22; mem['h0D9E]=8'h0A; mem['h0D9F]=8'h81;
    mem['h0DA0]=8'hD6; mem['h0DA1]=8'hAC; mem['h0DA2]=8'hD8; mem['h0DA3]=8'hFE;
    mem['h0DA4]=8'h07; mem['h0DA5]=8'hD0; mem['h0DA6]=8'h5F; mem['h0DA7]=8'h3A;
    mem['h0DA8]=8'hF2; mem['h0DA9]=8'h80; mem['h0DAA]=8'h3D; mem['h0DAB]=8'hB3;
    mem['h0DAC]=8'h7B; mem['h0DAD]=8'hCA; mem['h0DAE]=8'h1C; mem['h0DAF]=8'h13;
    mem['h0DB0]=8'h07; mem['h0DB1]=8'h83; mem['h0DB2]=8'h5F; mem['h0DB3]=8'h21;
    mem['h0DB4]=8'h7A; mem['h0DB5]=8'h03; mem['h0DB6]=8'h19; mem['h0DB7]=8'h78;
    mem['h0DB8]=8'h56; mem['h0DB9]=8'hBA; mem['h0DBA]=8'hD0; mem['h0DBB]=8'h23;
    mem['h0DBC]=8'hCD; mem['h0DBD]=8'h50; mem['h0DBE]=8'h0D; mem['h0DBF]=8'hC5;
    mem['h0DC0]=8'h01; mem['h0DC1]=8'h6E; mem['h0DC2]=8'h0D; mem['h0DC3]=8'hC5;
    mem['h0DC4]=8'h43; mem['h0DC5]=8'h4A; mem['h0DC6]=8'hCD; mem['h0DC7]=8'h60;
    mem['h0DC8]=8'h17; mem['h0DC9]=8'h58; mem['h0DCA]=8'h51; mem['h0DCB]=8'h4E;
    mem['h0DCC]=8'h23; mem['h0DCD]=8'h46; mem['h0DCE]=8'h23; mem['h0DCF]=8'hC5;
    mem['h0DD0]=8'h2A; mem['h0DD1]=8'h0A; mem['h0DD2]=8'h81; mem['h0DD3]=8'hC3;
    mem['h0DD4]=8'h62; mem['h0DD5]=8'h0D; mem['h0DD6]=8'hAF; mem['h0DD7]=8'h32;
    mem['h0DD8]=8'hF2; mem['h0DD9]=8'h80; mem['h0DDA]=8'hCD; mem['h0DDB]=8'hE0;
    mem['h0DDC]=8'h08; mem['h0DDD]=8'h1E; mem['h0DDE]=8'h24; mem['h0DDF]=8'hCA;
    mem['h0DE0]=8'h9C; mem['h0DE1]=8'h04; mem['h0DE2]=8'hDA; mem['h0DE3]=8'h36;
    mem['h0DE4]=8'h18; mem['h0DE5]=8'hCD; mem['h0DE6]=8'h7E; mem['h0DE7]=8'h09;
    mem['h0DE8]=8'hD2; mem['h0DE9]=8'h3D; mem['h0DEA]=8'h0E; mem['h0DEB]=8'hFE;
    mem['h0DEC]=8'h26; mem['h0DED]=8'h20; mem['h0DEE]=8'h12; mem['h0DEF]=8'hCD;
    mem['h0DF0]=8'hE0; mem['h0DF1]=8'h08; mem['h0DF2]=8'hFE; mem['h0DF3]=8'h48;
    mem['h0DF4]=8'hCA; mem['h0DF5]=8'h7A; mem['h0DF6]=8'h1C; mem['h0DF7]=8'hFE;
    mem['h0DF8]=8'h42; mem['h0DF9]=8'hCA; mem['h0DFA]=8'hEA; mem['h0DFB]=8'h1C;
    mem['h0DFC]=8'h1E; mem['h0DFD]=8'h02; mem['h0DFE]=8'hCA; mem['h0DFF]=8'h9C;
    mem['h0E00]=8'h04; mem['h0E01]=8'hFE; mem['h0E02]=8'hAC; mem['h0E03]=8'hCA;
    mem['h0E04]=8'hD6; mem['h0E05]=8'h0D; mem['h0E06]=8'hFE; mem['h0E07]=8'h2E;
    mem['h0E08]=8'hCA; mem['h0E09]=8'h36; mem['h0E0A]=8'h18; mem['h0E0B]=8'hFE;
    mem['h0E0C]=8'hAD; mem['h0E0D]=8'hCA; mem['h0E0E]=8'h2C; mem['h0E0F]=8'h0E;
    mem['h0E10]=8'hFE; mem['h0E11]=8'h22; mem['h0E12]=8'hCA; mem['h0E13]=8'hE5;
    mem['h0E14]=8'h11; mem['h0E15]=8'hFE; mem['h0E16]=8'hAA; mem['h0E17]=8'hCA;
    mem['h0E18]=8'h1E; mem['h0E19]=8'h0F; mem['h0E1A]=8'hFE; mem['h0E1B]=8'hA7;
    mem['h0E1C]=8'hCA; mem['h0E1D]=8'h49; mem['h0E1E]=8'h11; mem['h0E1F]=8'hD6;
    mem['h0E20]=8'hB6; mem['h0E21]=8'hD2; mem['h0E22]=8'h4E; mem['h0E23]=8'h0E;
    mem['h0E24]=8'hCD; mem['h0E25]=8'h5B; mem['h0E26]=8'h0D; mem['h0E27]=8'hCD;
    mem['h0E28]=8'h56; mem['h0E29]=8'h07; mem['h0E2A]=8'h29; mem['h0E2B]=8'hC9;
    mem['h0E2C]=8'h16; mem['h0E2D]=8'h7D; mem['h0E2E]=8'hCD; mem['h0E2F]=8'h62;
    mem['h0E30]=8'h0D; mem['h0E31]=8'h2A; mem['h0E32]=8'h15; mem['h0E33]=8'h81;
    mem['h0E34]=8'hE5; mem['h0E35]=8'hCD; mem['h0E36]=8'h58; mem['h0E37]=8'h17;
    mem['h0E38]=8'hCD; mem['h0E39]=8'h50; mem['h0E3A]=8'h0D; mem['h0E3B]=8'hE1;
    mem['h0E3C]=8'hC9; mem['h0E3D]=8'hCD; mem['h0E3E]=8'h43; mem['h0E3F]=8'h0F;
    mem['h0E40]=8'hE5; mem['h0E41]=8'hEB; mem['h0E42]=8'h22; mem['h0E43]=8'h29;
    mem['h0E44]=8'h81; mem['h0E45]=8'h3A; mem['h0E46]=8'hF2; mem['h0E47]=8'h80;
    mem['h0E48]=8'hB7; mem['h0E49]=8'hCC; mem['h0E4A]=8'h6D; mem['h0E4B]=8'h17;
    mem['h0E4C]=8'hE1; mem['h0E4D]=8'hC9; mem['h0E4E]=8'h06; mem['h0E4F]=8'h00;
    mem['h0E50]=8'h07; mem['h0E51]=8'h4F; mem['h0E52]=8'hC5; mem['h0E53]=8'hCD;
    mem['h0E54]=8'hE0; mem['h0E55]=8'h08; mem['h0E56]=8'h79; mem['h0E57]=8'hFE;
    mem['h0E58]=8'h31; mem['h0E59]=8'hDA; mem['h0E5A]=8'h75; mem['h0E5B]=8'h0E;
    mem['h0E5C]=8'hCD; mem['h0E5D]=8'h5B; mem['h0E5E]=8'h0D; mem['h0E5F]=8'hCD;
    mem['h0E60]=8'h56; mem['h0E61]=8'h07; mem['h0E62]=8'h2C; mem['h0E63]=8'hCD;
    mem['h0E64]=8'h51; mem['h0E65]=8'h0D; mem['h0E66]=8'hEB; mem['h0E67]=8'h2A;
    mem['h0E68]=8'h29; mem['h0E69]=8'h81; mem['h0E6A]=8'hE3; mem['h0E6B]=8'hE5;
    mem['h0E6C]=8'hEB; mem['h0E6D]=8'hCD; mem['h0E6E]=8'hAE; mem['h0E6F]=8'h14;
    mem['h0E70]=8'hEB; mem['h0E71]=8'hE3; mem['h0E72]=8'hC3; mem['h0E73]=8'h7D;
    mem['h0E74]=8'h0E; mem['h0E75]=8'hCD; mem['h0E76]=8'h24; mem['h0E77]=8'h0E;
    mem['h0E78]=8'hE3; mem['h0E79]=8'h11; mem['h0E7A]=8'h38; mem['h0E7B]=8'h0E;
    mem['h0E7C]=8'hD5; mem['h0E7D]=8'h01; mem['h0E7E]=8'hD9; mem['h0E7F]=8'h01;
    mem['h0E80]=8'h09; mem['h0E81]=8'h4E; mem['h0E82]=8'h23; mem['h0E83]=8'h66;
    mem['h0E84]=8'h69; mem['h0E85]=8'hE9; mem['h0E86]=8'h15; mem['h0E87]=8'hFE;
    mem['h0E88]=8'hAD; mem['h0E89]=8'hC8; mem['h0E8A]=8'hFE; mem['h0E8B]=8'h2D;
    mem['h0E8C]=8'hC8; mem['h0E8D]=8'h14; mem['h0E8E]=8'hFE; mem['h0E8F]=8'h2B;
    mem['h0E90]=8'hC8; mem['h0E91]=8'hFE; mem['h0E92]=8'hAC; mem['h0E93]=8'hC8;
    mem['h0E94]=8'h2B; mem['h0E95]=8'hC9; mem['h0E96]=8'hF6; mem['h0E97]=8'hAF;
    mem['h0E98]=8'hF5; mem['h0E99]=8'hCD; mem['h0E9A]=8'h50; mem['h0E9B]=8'h0D;
    mem['h0E9C]=8'hCD; mem['h0E9D]=8'h92; mem['h0E9E]=8'h09; mem['h0E9F]=8'hF1;
    mem['h0EA0]=8'hEB; mem['h0EA1]=8'hC1; mem['h0EA2]=8'hE3; mem['h0EA3]=8'hEB;
    mem['h0EA4]=8'hCD; mem['h0EA5]=8'h70; mem['h0EA6]=8'h17; mem['h0EA7]=8'hF5;
    mem['h0EA8]=8'hCD; mem['h0EA9]=8'h92; mem['h0EAA]=8'h09; mem['h0EAB]=8'hF1;
    mem['h0EAC]=8'hC1; mem['h0EAD]=8'h79; mem['h0EAE]=8'h21; mem['h0EAF]=8'h07;
    mem['h0EB0]=8'h11; mem['h0EB1]=8'hC2; mem['h0EB2]=8'hB9; mem['h0EB3]=8'h0E;
    mem['h0EB4]=8'hA3; mem['h0EB5]=8'h4F; mem['h0EB6]=8'h78; mem['h0EB7]=8'hA2;
    mem['h0EB8]=8'hE9; mem['h0EB9]=8'hB3; mem['h0EBA]=8'h4F; mem['h0EBB]=8'h78;
    mem['h0EBC]=8'hB2; mem['h0EBD]=8'hE9; mem['h0EBE]=8'h21; mem['h0EBF]=8'hD0;
    mem['h0EC0]=8'h0E; mem['h0EC1]=8'h3A; mem['h0EC2]=8'hF2; mem['h0EC3]=8'h80;
    mem['h0EC4]=8'h1F; mem['h0EC5]=8'h7A; mem['h0EC6]=8'h17; mem['h0EC7]=8'h5F;
    mem['h0EC8]=8'h16; mem['h0EC9]=8'h64; mem['h0ECA]=8'h78; mem['h0ECB]=8'hBA;
    mem['h0ECC]=8'hD0; mem['h0ECD]=8'hC3; mem['h0ECE]=8'hBF; mem['h0ECF]=8'h0D;
    mem['h0ED0]=8'hD2; mem['h0ED1]=8'h0E; mem['h0ED2]=8'h79; mem['h0ED3]=8'hB7;
    mem['h0ED4]=8'h1F; mem['h0ED5]=8'hC1; mem['h0ED6]=8'hD1; mem['h0ED7]=8'hF5;
    mem['h0ED8]=8'hCD; mem['h0ED9]=8'h52; mem['h0EDA]=8'h0D; mem['h0EDB]=8'h21;
    mem['h0EDC]=8'h14; mem['h0EDD]=8'h0F; mem['h0EDE]=8'hE5; mem['h0EDF]=8'hCA;
    mem['h0EE0]=8'hAA; mem['h0EE1]=8'h17; mem['h0EE2]=8'hAF; mem['h0EE3]=8'h32;
    mem['h0EE4]=8'hF2; mem['h0EE5]=8'h80; mem['h0EE6]=8'hD5; mem['h0EE7]=8'hCD;
    mem['h0EE8]=8'h69; mem['h0EE9]=8'h13; mem['h0EEA]=8'h7E; mem['h0EEB]=8'h23;
    mem['h0EEC]=8'h23; mem['h0EED]=8'h4E; mem['h0EEE]=8'h23; mem['h0EEF]=8'h46;
    mem['h0EF0]=8'hD1; mem['h0EF1]=8'hC5; mem['h0EF2]=8'hF5; mem['h0EF3]=8'hCD;
    mem['h0EF4]=8'h6D; mem['h0EF5]=8'h13; mem['h0EF6]=8'hCD; mem['h0EF7]=8'h7E;
    mem['h0EF8]=8'h17; mem['h0EF9]=8'hF1; mem['h0EFA]=8'h57; mem['h0EFB]=8'hE1;
    mem['h0EFC]=8'h7B; mem['h0EFD]=8'hB2; mem['h0EFE]=8'hC8; mem['h0EFF]=8'h7A;
    mem['h0F00]=8'hD6; mem['h0F01]=8'h01; mem['h0F02]=8'hD8; mem['h0F03]=8'hAF;
    mem['h0F04]=8'hBB; mem['h0F05]=8'h3C; mem['h0F06]=8'hD0; mem['h0F07]=8'h15;
    mem['h0F08]=8'h1D; mem['h0F09]=8'h0A; mem['h0F0A]=8'hBE; mem['h0F0B]=8'h23;
    mem['h0F0C]=8'h03; mem['h0F0D]=8'hCA; mem['h0F0E]=8'hFC; mem['h0F0F]=8'h0E;
    mem['h0F10]=8'h3F; mem['h0F11]=8'hC3; mem['h0F12]=8'h3A; mem['h0F13]=8'h17;
    mem['h0F14]=8'h3C; mem['h0F15]=8'h8F; mem['h0F16]=8'hC1; mem['h0F17]=8'hA0;
    mem['h0F18]=8'hC6; mem['h0F19]=8'hFF; mem['h0F1A]=8'h9F; mem['h0F1B]=8'hC3;
    mem['h0F1C]=8'h41; mem['h0F1D]=8'h17; mem['h0F1E]=8'h16; mem['h0F1F]=8'h5A;
    mem['h0F20]=8'hCD; mem['h0F21]=8'h62; mem['h0F22]=8'h0D; mem['h0F23]=8'hCD;
    mem['h0F24]=8'h50; mem['h0F25]=8'h0D; mem['h0F26]=8'hCD; mem['h0F27]=8'h92;
    mem['h0F28]=8'h09; mem['h0F29]=8'h7B; mem['h0F2A]=8'h2F; mem['h0F2B]=8'h4F;
    mem['h0F2C]=8'h7A; mem['h0F2D]=8'h2F; mem['h0F2E]=8'hCD; mem['h0F2F]=8'h07;
    mem['h0F30]=8'h11; mem['h0F31]=8'hC1; mem['h0F32]=8'hC3; mem['h0F33]=8'h6E;
    mem['h0F34]=8'h0D; mem['h0F35]=8'h2B; mem['h0F36]=8'hCD; mem['h0F37]=8'hE0;
    mem['h0F38]=8'h08; mem['h0F39]=8'hC8; mem['h0F3A]=8'hCD; mem['h0F3B]=8'h56;
    mem['h0F3C]=8'h07; mem['h0F3D]=8'h2C; mem['h0F3E]=8'h01; mem['h0F3F]=8'h35;
    mem['h0F40]=8'h0F; mem['h0F41]=8'hC5; mem['h0F42]=8'hF6; mem['h0F43]=8'hAF;
    mem['h0F44]=8'h32; mem['h0F45]=8'hF1; mem['h0F46]=8'h80; mem['h0F47]=8'h46;
    mem['h0F48]=8'hCD; mem['h0F49]=8'h7E; mem['h0F4A]=8'h09; mem['h0F4B]=8'hDA;
    mem['h0F4C]=8'h88; mem['h0F4D]=8'h04; mem['h0F4E]=8'hAF; mem['h0F4F]=8'h4F;
    mem['h0F50]=8'h32; mem['h0F51]=8'hF2; mem['h0F52]=8'h80; mem['h0F53]=8'hCD;
    mem['h0F54]=8'hE0; mem['h0F55]=8'h08; mem['h0F56]=8'hDA; mem['h0F57]=8'h5F;
    mem['h0F58]=8'h0F; mem['h0F59]=8'hCD; mem['h0F5A]=8'h7E; mem['h0F5B]=8'h09;
    mem['h0F5C]=8'hDA; mem['h0F5D]=8'h6C; mem['h0F5E]=8'h0F; mem['h0F5F]=8'h4F;
    mem['h0F60]=8'hCD; mem['h0F61]=8'hE0; mem['h0F62]=8'h08; mem['h0F63]=8'hDA;
    mem['h0F64]=8'h60; mem['h0F65]=8'h0F; mem['h0F66]=8'hCD; mem['h0F67]=8'h7E;
    mem['h0F68]=8'h09; mem['h0F69]=8'hD2; mem['h0F6A]=8'h60; mem['h0F6B]=8'h0F;
    mem['h0F6C]=8'hD6; mem['h0F6D]=8'h24; mem['h0F6E]=8'hC2; mem['h0F6F]=8'h7B;
    mem['h0F70]=8'h0F; mem['h0F71]=8'h3C; mem['h0F72]=8'h32; mem['h0F73]=8'hF2;
    mem['h0F74]=8'h80; mem['h0F75]=8'h0F; mem['h0F76]=8'h81; mem['h0F77]=8'h4F;
    mem['h0F78]=8'hCD; mem['h0F79]=8'hE0; mem['h0F7A]=8'h08; mem['h0F7B]=8'h3A;
    mem['h0F7C]=8'h10; mem['h0F7D]=8'h81; mem['h0F7E]=8'h3D; mem['h0F7F]=8'hCA;
    mem['h0F80]=8'h28; mem['h0F81]=8'h10; mem['h0F82]=8'hF2; mem['h0F83]=8'h8B;
    mem['h0F84]=8'h0F; mem['h0F85]=8'h7E; mem['h0F86]=8'hD6; mem['h0F87]=8'h28;
    mem['h0F88]=8'hCA; mem['h0F89]=8'h00; mem['h0F8A]=8'h10; mem['h0F8B]=8'hAF;
    mem['h0F8C]=8'h32; mem['h0F8D]=8'h10; mem['h0F8E]=8'h81; mem['h0F8F]=8'hE5;
    mem['h0F90]=8'h50; mem['h0F91]=8'h59; mem['h0F92]=8'h2A; mem['h0F93]=8'h23;
    mem['h0F94]=8'h81; mem['h0F95]=8'hCD; mem['h0F96]=8'h50; mem['h0F97]=8'h07;
    mem['h0F98]=8'h11; mem['h0F99]=8'h25; mem['h0F9A]=8'h81; mem['h0F9B]=8'hCA;
    mem['h0F9C]=8'h70; mem['h0F9D]=8'h16; mem['h0F9E]=8'h2A; mem['h0F9F]=8'h1D;
    mem['h0FA0]=8'h81; mem['h0FA1]=8'hEB; mem['h0FA2]=8'h2A; mem['h0FA3]=8'h1B;
    mem['h0FA4]=8'h81; mem['h0FA5]=8'hCD; mem['h0FA6]=8'h50; mem['h0FA7]=8'h07;
    mem['h0FA8]=8'hCA; mem['h0FA9]=8'hBE; mem['h0FAA]=8'h0F; mem['h0FAB]=8'h79;
    mem['h0FAC]=8'h96; mem['h0FAD]=8'h23; mem['h0FAE]=8'hC2; mem['h0FAF]=8'hB3;
    mem['h0FB0]=8'h0F; mem['h0FB1]=8'h78; mem['h0FB2]=8'h96; mem['h0FB3]=8'h23;
    mem['h0FB4]=8'hCA; mem['h0FB5]=8'hF2; mem['h0FB6]=8'h0F; mem['h0FB7]=8'h23;
    mem['h0FB8]=8'h23; mem['h0FB9]=8'h23; mem['h0FBA]=8'h23; mem['h0FBB]=8'hC3;
    mem['h0FBC]=8'hA5; mem['h0FBD]=8'h0F; mem['h0FBE]=8'hE1; mem['h0FBF]=8'hE3;
    mem['h0FC0]=8'hD5; mem['h0FC1]=8'h11; mem['h0FC2]=8'h40; mem['h0FC3]=8'h0E;
    mem['h0FC4]=8'hCD; mem['h0FC5]=8'h50; mem['h0FC6]=8'h07; mem['h0FC7]=8'hD1;
    mem['h0FC8]=8'hCA; mem['h0FC9]=8'hF5; mem['h0FCA]=8'h0F; mem['h0FCB]=8'hE3;
    mem['h0FCC]=8'hE5; mem['h0FCD]=8'hC5; mem['h0FCE]=8'h01; mem['h0FCF]=8'h06;
    mem['h0FD0]=8'h00; mem['h0FD1]=8'h2A; mem['h0FD2]=8'h1F; mem['h0FD3]=8'h81;
    mem['h0FD4]=8'hE5; mem['h0FD5]=8'h09; mem['h0FD6]=8'hC1; mem['h0FD7]=8'hE5;
    mem['h0FD8]=8'hCD; mem['h0FD9]=8'h54; mem['h0FDA]=8'h04; mem['h0FDB]=8'hE1;
    mem['h0FDC]=8'h22; mem['h0FDD]=8'h1F; mem['h0FDE]=8'h81; mem['h0FDF]=8'h60;
    mem['h0FE0]=8'h69; mem['h0FE1]=8'h22; mem['h0FE2]=8'h1D; mem['h0FE3]=8'h81;
    mem['h0FE4]=8'h2B; mem['h0FE5]=8'h36; mem['h0FE6]=8'h00; mem['h0FE7]=8'hCD;
    mem['h0FE8]=8'h50; mem['h0FE9]=8'h07; mem['h0FEA]=8'hC2; mem['h0FEB]=8'hE4;
    mem['h0FEC]=8'h0F; mem['h0FED]=8'hD1; mem['h0FEE]=8'h73; mem['h0FEF]=8'h23;
    mem['h0FF0]=8'h72; mem['h0FF1]=8'h23; mem['h0FF2]=8'hEB; mem['h0FF3]=8'hE1;
    mem['h0FF4]=8'hC9; mem['h0FF5]=8'h32; mem['h0FF6]=8'h2C; mem['h0FF7]=8'h81;
    mem['h0FF8]=8'h21; mem['h0FF9]=8'h24; mem['h0FFA]=8'h04; mem['h0FFB]=8'h22;
    mem['h0FFC]=8'h29; mem['h0FFD]=8'h81; mem['h0FFE]=8'hE1; mem['h0FFF]=8'hC9;
    mem['h1000]=8'hE5; mem['h1001]=8'h2A; mem['h1002]=8'hF1; mem['h1003]=8'h80;
    mem['h1004]=8'hE3; mem['h1005]=8'h57; mem['h1006]=8'hD5; mem['h1007]=8'hC5;
    mem['h1008]=8'hCD; mem['h1009]=8'h86; mem['h100A]=8'h09; mem['h100B]=8'hC1;
    mem['h100C]=8'hF1; mem['h100D]=8'hEB; mem['h100E]=8'hE3; mem['h100F]=8'hE5;
    mem['h1010]=8'hEB; mem['h1011]=8'h3C; mem['h1012]=8'h57; mem['h1013]=8'h7E;
    mem['h1014]=8'hFE; mem['h1015]=8'h2C; mem['h1016]=8'hCA; mem['h1017]=8'h06;
    mem['h1018]=8'h10; mem['h1019]=8'hCD; mem['h101A]=8'h56; mem['h101B]=8'h07;
    mem['h101C]=8'h29; mem['h101D]=8'h22; mem['h101E]=8'h15; mem['h101F]=8'h81;
    mem['h1020]=8'hE1; mem['h1021]=8'h22; mem['h1022]=8'hF1; mem['h1023]=8'h80;
    mem['h1024]=8'h1E; mem['h1025]=8'h00; mem['h1026]=8'hD5; mem['h1027]=8'h11;
    mem['h1028]=8'hE5; mem['h1029]=8'hF5; mem['h102A]=8'h2A; mem['h102B]=8'h1D;
    mem['h102C]=8'h81; mem['h102D]=8'h3E; mem['h102E]=8'h19; mem['h102F]=8'hEB;
    mem['h1030]=8'h2A; mem['h1031]=8'h1F; mem['h1032]=8'h81; mem['h1033]=8'hEB;
    mem['h1034]=8'hCD; mem['h1035]=8'h50; mem['h1036]=8'h07; mem['h1037]=8'hCA;
    mem['h1038]=8'h60; mem['h1039]=8'h10; mem['h103A]=8'h7E; mem['h103B]=8'hB9;
    mem['h103C]=8'h23; mem['h103D]=8'hC2; mem['h103E]=8'h42; mem['h103F]=8'h10;
    mem['h1040]=8'h7E; mem['h1041]=8'hB8; mem['h1042]=8'h23; mem['h1043]=8'h5E;
    mem['h1044]=8'h23; mem['h1045]=8'h56; mem['h1046]=8'h23; mem['h1047]=8'hC2;
    mem['h1048]=8'h2E; mem['h1049]=8'h10; mem['h104A]=8'h3A; mem['h104B]=8'hF1;
    mem['h104C]=8'h80; mem['h104D]=8'hB7; mem['h104E]=8'hC2; mem['h104F]=8'h91;
    mem['h1050]=8'h04; mem['h1051]=8'hF1; mem['h1052]=8'h44; mem['h1053]=8'h4D;
    mem['h1054]=8'hCA; mem['h1055]=8'h70; mem['h1056]=8'h16; mem['h1057]=8'h96;
    mem['h1058]=8'hCA; mem['h1059]=8'hBE; mem['h105A]=8'h10; mem['h105B]=8'h1E;
    mem['h105C]=8'h10; mem['h105D]=8'hC3; mem['h105E]=8'h9C; mem['h105F]=8'h04;
    mem['h1060]=8'h11; mem['h1061]=8'h04; mem['h1062]=8'h00; mem['h1063]=8'hF1;
    mem['h1064]=8'hCA; mem['h1065]=8'hA7; mem['h1066]=8'h09; mem['h1067]=8'h71;
    mem['h1068]=8'h23; mem['h1069]=8'h70; mem['h106A]=8'h23; mem['h106B]=8'h4F;
    mem['h106C]=8'hCD; mem['h106D]=8'h65; mem['h106E]=8'h04; mem['h106F]=8'h23;
    mem['h1070]=8'h23; mem['h1071]=8'h22; mem['h1072]=8'h0A; mem['h1073]=8'h81;
    mem['h1074]=8'h71; mem['h1075]=8'h23; mem['h1076]=8'h3A; mem['h1077]=8'hF1;
    mem['h1078]=8'h80; mem['h1079]=8'h17; mem['h107A]=8'h79; mem['h107B]=8'h01;
    mem['h107C]=8'h0B; mem['h107D]=8'h00; mem['h107E]=8'hD2; mem['h107F]=8'h83;
    mem['h1080]=8'h10; mem['h1081]=8'hC1; mem['h1082]=8'h03; mem['h1083]=8'h71;
    mem['h1084]=8'h23; mem['h1085]=8'h70; mem['h1086]=8'h23; mem['h1087]=8'hF5;
    mem['h1088]=8'hE5; mem['h1089]=8'hCD; mem['h108A]=8'h1B; mem['h108B]=8'h18;
    mem['h108C]=8'hEB; mem['h108D]=8'hE1; mem['h108E]=8'hF1; mem['h108F]=8'h3D;
    mem['h1090]=8'hC2; mem['h1091]=8'h7B; mem['h1092]=8'h10; mem['h1093]=8'hF5;
    mem['h1094]=8'h42; mem['h1095]=8'h4B; mem['h1096]=8'hEB; mem['h1097]=8'h19;
    mem['h1098]=8'hDA; mem['h1099]=8'h7D; mem['h109A]=8'h04; mem['h109B]=8'hCD;
    mem['h109C]=8'h6E; mem['h109D]=8'h04; mem['h109E]=8'h22; mem['h109F]=8'h1F;
    mem['h10A0]=8'h81; mem['h10A1]=8'h2B; mem['h10A2]=8'h36; mem['h10A3]=8'h00;
    mem['h10A4]=8'hCD; mem['h10A5]=8'h50; mem['h10A6]=8'h07; mem['h10A7]=8'hC2;
    mem['h10A8]=8'hA1; mem['h10A9]=8'h10; mem['h10AA]=8'h03; mem['h10AB]=8'h57;
    mem['h10AC]=8'h2A; mem['h10AD]=8'h0A; mem['h10AE]=8'h81; mem['h10AF]=8'h5E;
    mem['h10B0]=8'hEB; mem['h10B1]=8'h29; mem['h10B2]=8'h09; mem['h10B3]=8'hEB;
    mem['h10B4]=8'h2B; mem['h10B5]=8'h2B; mem['h10B6]=8'h73; mem['h10B7]=8'h23;
    mem['h10B8]=8'h72; mem['h10B9]=8'h23; mem['h10BA]=8'hF1; mem['h10BB]=8'hDA;
    mem['h10BC]=8'hE2; mem['h10BD]=8'h10; mem['h10BE]=8'h47; mem['h10BF]=8'h4F;
    mem['h10C0]=8'h7E; mem['h10C1]=8'h23; mem['h10C2]=8'h16; mem['h10C3]=8'hE1;
    mem['h10C4]=8'h5E; mem['h10C5]=8'h23; mem['h10C6]=8'h56; mem['h10C7]=8'h23;
    mem['h10C8]=8'hE3; mem['h10C9]=8'hF5; mem['h10CA]=8'hCD; mem['h10CB]=8'h50;
    mem['h10CC]=8'h07; mem['h10CD]=8'hD2; mem['h10CE]=8'h5B; mem['h10CF]=8'h10;
    mem['h10D0]=8'hE5; mem['h10D1]=8'hCD; mem['h10D2]=8'h1B; mem['h10D3]=8'h18;
    mem['h10D4]=8'hD1; mem['h10D5]=8'h19; mem['h10D6]=8'hF1; mem['h10D7]=8'h3D;
    mem['h10D8]=8'h44; mem['h10D9]=8'h4D; mem['h10DA]=8'hC2; mem['h10DB]=8'hC3;
    mem['h10DC]=8'h10; mem['h10DD]=8'h29; mem['h10DE]=8'h29; mem['h10DF]=8'hC1;
    mem['h10E0]=8'h09; mem['h10E1]=8'hEB; mem['h10E2]=8'h2A; mem['h10E3]=8'h15;
    mem['h10E4]=8'h81; mem['h10E5]=8'hC9; mem['h10E6]=8'h2A; mem['h10E7]=8'h1F;
    mem['h10E8]=8'h81; mem['h10E9]=8'hEB; mem['h10EA]=8'h21; mem['h10EB]=8'h00;
    mem['h10EC]=8'h00; mem['h10ED]=8'h39; mem['h10EE]=8'h3A; mem['h10EF]=8'hF2;
    mem['h10F0]=8'h80; mem['h10F1]=8'hB7; mem['h10F2]=8'hCA; mem['h10F3]=8'h02;
    mem['h10F4]=8'h11; mem['h10F5]=8'hCD; mem['h10F6]=8'h69; mem['h10F7]=8'h13;
    mem['h10F8]=8'hCD; mem['h10F9]=8'h69; mem['h10FA]=8'h12; mem['h10FB]=8'h2A;
    mem['h10FC]=8'h9F; mem['h10FD]=8'h80; mem['h10FE]=8'hEB; mem['h10FF]=8'h2A;
    mem['h1100]=8'h08; mem['h1101]=8'h81; mem['h1102]=8'h7D; mem['h1103]=8'h93;
    mem['h1104]=8'h4F; mem['h1105]=8'h7C; mem['h1106]=8'h9A; mem['h1107]=8'h41;
    mem['h1108]=8'h50; mem['h1109]=8'h1E; mem['h110A]=8'h00; mem['h110B]=8'h21;
    mem['h110C]=8'hF2; mem['h110D]=8'h80; mem['h110E]=8'h73; mem['h110F]=8'h06;
    mem['h1110]=8'h90; mem['h1111]=8'hC3; mem['h1112]=8'h46; mem['h1113]=8'h17;
    mem['h1114]=8'h3A; mem['h1115]=8'hF0; mem['h1116]=8'h80; mem['h1117]=8'h47;
    mem['h1118]=8'hAF; mem['h1119]=8'hC3; mem['h111A]=8'h08; mem['h111B]=8'h11;
    mem['h111C]=8'hCD; mem['h111D]=8'h9F; mem['h111E]=8'h11; mem['h111F]=8'hCD;
    mem['h1120]=8'h91; mem['h1121]=8'h11; mem['h1122]=8'h01; mem['h1123]=8'h77;
    mem['h1124]=8'h0A; mem['h1125]=8'hC5; mem['h1126]=8'hD5; mem['h1127]=8'hCD;
    mem['h1128]=8'h56; mem['h1129]=8'h07; mem['h112A]=8'h28; mem['h112B]=8'hCD;
    mem['h112C]=8'h43; mem['h112D]=8'h0F; mem['h112E]=8'hE5; mem['h112F]=8'hEB;
    mem['h1130]=8'h2B; mem['h1131]=8'h56; mem['h1132]=8'h2B; mem['h1133]=8'h5E;
    mem['h1134]=8'hE1; mem['h1135]=8'hCD; mem['h1136]=8'h50; mem['h1137]=8'h0D;
    mem['h1138]=8'hCD; mem['h1139]=8'h56; mem['h113A]=8'h07; mem['h113B]=8'h29;
    mem['h113C]=8'hCD; mem['h113D]=8'h56; mem['h113E]=8'h07; mem['h113F]=8'hB4;
    mem['h1140]=8'h44; mem['h1141]=8'h4D; mem['h1142]=8'hE3; mem['h1143]=8'h71;
    mem['h1144]=8'h23; mem['h1145]=8'h70; mem['h1146]=8'hC3; mem['h1147]=8'hDE;
    mem['h1148]=8'h11; mem['h1149]=8'hCD; mem['h114A]=8'h9F; mem['h114B]=8'h11;
    mem['h114C]=8'hD5; mem['h114D]=8'hCD; mem['h114E]=8'h24; mem['h114F]=8'h0E;
    mem['h1150]=8'hCD; mem['h1151]=8'h50; mem['h1152]=8'h0D; mem['h1153]=8'hE3;
    mem['h1154]=8'h5E; mem['h1155]=8'h23; mem['h1156]=8'h56; mem['h1157]=8'h23;
    mem['h1158]=8'h7A; mem['h1159]=8'hB3; mem['h115A]=8'hCA; mem['h115B]=8'h94;
    mem['h115C]=8'h04; mem['h115D]=8'h7E; mem['h115E]=8'h23; mem['h115F]=8'h66;
    mem['h1160]=8'h6F; mem['h1161]=8'hE5; mem['h1162]=8'h2A; mem['h1163]=8'h23;
    mem['h1164]=8'h81; mem['h1165]=8'hE3; mem['h1166]=8'h22; mem['h1167]=8'h23;
    mem['h1168]=8'h81; mem['h1169]=8'h2A; mem['h116A]=8'h27; mem['h116B]=8'h81;
    mem['h116C]=8'hE5; mem['h116D]=8'h2A; mem['h116E]=8'h25; mem['h116F]=8'h81;
    mem['h1170]=8'hE5; mem['h1171]=8'h21; mem['h1172]=8'h25; mem['h1173]=8'h81;
    mem['h1174]=8'hD5; mem['h1175]=8'hCD; mem['h1176]=8'h87; mem['h1177]=8'h17;
    mem['h1178]=8'hE1; mem['h1179]=8'hCD; mem['h117A]=8'h4D; mem['h117B]=8'h0D;
    mem['h117C]=8'h2B; mem['h117D]=8'hCD; mem['h117E]=8'hE0; mem['h117F]=8'h08;
    mem['h1180]=8'hC2; mem['h1181]=8'h88; mem['h1182]=8'h04; mem['h1183]=8'hE1;
    mem['h1184]=8'h22; mem['h1185]=8'h25; mem['h1186]=8'h81; mem['h1187]=8'hE1;
    mem['h1188]=8'h22; mem['h1189]=8'h27; mem['h118A]=8'h81; mem['h118B]=8'hE1;
    mem['h118C]=8'h22; mem['h118D]=8'h23; mem['h118E]=8'h81; mem['h118F]=8'hE1;
    mem['h1190]=8'hC9; mem['h1191]=8'hE5; mem['h1192]=8'h2A; mem['h1193]=8'hA1;
    mem['h1194]=8'h80; mem['h1195]=8'h23; mem['h1196]=8'h7C; mem['h1197]=8'hB5;
    mem['h1198]=8'hE1; mem['h1199]=8'hC0; mem['h119A]=8'h1E; mem['h119B]=8'h16;
    mem['h119C]=8'hC3; mem['h119D]=8'h9C; mem['h119E]=8'h04; mem['h119F]=8'hCD;
    mem['h11A0]=8'h56; mem['h11A1]=8'h07; mem['h11A2]=8'hA7; mem['h11A3]=8'h3E;
    mem['h11A4]=8'h80; mem['h11A5]=8'h32; mem['h11A6]=8'h10; mem['h11A7]=8'h81;
    mem['h11A8]=8'hB6; mem['h11A9]=8'h47; mem['h11AA]=8'hCD; mem['h11AB]=8'h48;
    mem['h11AC]=8'h0F; mem['h11AD]=8'hC3; mem['h11AE]=8'h50; mem['h11AF]=8'h0D;
    mem['h11B0]=8'hCD; mem['h11B1]=8'h50; mem['h11B2]=8'h0D; mem['h11B3]=8'hCD;
    mem['h11B4]=8'hD4; mem['h11B5]=8'h18; mem['h11B6]=8'hCD; mem['h11B7]=8'hE4;
    mem['h11B8]=8'h11; mem['h11B9]=8'hCD; mem['h11BA]=8'h69; mem['h11BB]=8'h13;
    mem['h11BC]=8'h01; mem['h11BD]=8'hC4; mem['h11BE]=8'h13; mem['h11BF]=8'hC5;
    mem['h11C0]=8'h7E; mem['h11C1]=8'h23; mem['h11C2]=8'h23; mem['h11C3]=8'hE5;
    mem['h11C4]=8'hCD; mem['h11C5]=8'h3F; mem['h11C6]=8'h12; mem['h11C7]=8'hE1;
    mem['h11C8]=8'h4E; mem['h11C9]=8'h23; mem['h11CA]=8'h46; mem['h11CB]=8'hCD;
    mem['h11CC]=8'hD8; mem['h11CD]=8'h11; mem['h11CE]=8'hE5; mem['h11CF]=8'h6F;
    mem['h11D0]=8'hCD; mem['h11D1]=8'h5C; mem['h11D2]=8'h13; mem['h11D3]=8'hD1;
    mem['h11D4]=8'hC9; mem['h11D5]=8'hCD; mem['h11D6]=8'h3F; mem['h11D7]=8'h12;
    mem['h11D8]=8'h21; mem['h11D9]=8'h04; mem['h11DA]=8'h81; mem['h11DB]=8'hE5;
    mem['h11DC]=8'h77; mem['h11DD]=8'h23; mem['h11DE]=8'h23; mem['h11DF]=8'h73;
    mem['h11E0]=8'h23; mem['h11E1]=8'h72; mem['h11E2]=8'hE1; mem['h11E3]=8'hC9;
    mem['h11E4]=8'h2B; mem['h11E5]=8'h06; mem['h11E6]=8'h22; mem['h11E7]=8'h50;
    mem['h11E8]=8'hE5; mem['h11E9]=8'h0E; mem['h11EA]=8'hFF; mem['h11EB]=8'h23;
    mem['h11EC]=8'h7E; mem['h11ED]=8'h0C; mem['h11EE]=8'hB7; mem['h11EF]=8'hCA;
    mem['h11F0]=8'hFA; mem['h11F1]=8'h11; mem['h11F2]=8'hBA; mem['h11F3]=8'hCA;
    mem['h11F4]=8'hFA; mem['h11F5]=8'h11; mem['h11F6]=8'hB8; mem['h11F7]=8'hC2;
    mem['h11F8]=8'hEB; mem['h11F9]=8'h11; mem['h11FA]=8'hFE; mem['h11FB]=8'h22;
    mem['h11FC]=8'hCC; mem['h11FD]=8'hE0; mem['h11FE]=8'h08; mem['h11FF]=8'hE3;
    mem['h1200]=8'h23; mem['h1201]=8'hEB; mem['h1202]=8'h79; mem['h1203]=8'hCD;
    mem['h1204]=8'hD8; mem['h1205]=8'h11; mem['h1206]=8'h11; mem['h1207]=8'h04;
    mem['h1208]=8'h81; mem['h1209]=8'h2A; mem['h120A]=8'hF6; mem['h120B]=8'h80;
    mem['h120C]=8'h22; mem['h120D]=8'h29; mem['h120E]=8'h81; mem['h120F]=8'h3E;
    mem['h1210]=8'h01; mem['h1211]=8'h32; mem['h1212]=8'hF2; mem['h1213]=8'h80;
    mem['h1214]=8'hCD; mem['h1215]=8'h8A; mem['h1216]=8'h17; mem['h1217]=8'hCD;
    mem['h1218]=8'h50; mem['h1219]=8'h07; mem['h121A]=8'h22; mem['h121B]=8'hF6;
    mem['h121C]=8'h80; mem['h121D]=8'hE1; mem['h121E]=8'h7E; mem['h121F]=8'hC0;
    mem['h1220]=8'h1E; mem['h1221]=8'h1E; mem['h1222]=8'hC3; mem['h1223]=8'h9C;
    mem['h1224]=8'h04; mem['h1225]=8'h23; mem['h1226]=8'hCD; mem['h1227]=8'hE4;
    mem['h1228]=8'h11; mem['h1229]=8'hCD; mem['h122A]=8'h69; mem['h122B]=8'h13;
    mem['h122C]=8'hCD; mem['h122D]=8'h7E; mem['h122E]=8'h17; mem['h122F]=8'h1C;
    mem['h1230]=8'h1D; mem['h1231]=8'hC8; mem['h1232]=8'h0A; mem['h1233]=8'hCD;
    mem['h1234]=8'h61; mem['h1235]=8'h07; mem['h1236]=8'hFE; mem['h1237]=8'h0D;
    mem['h1238]=8'hCC; mem['h1239]=8'h92; mem['h123A]=8'h0B; mem['h123B]=8'h03;
    mem['h123C]=8'hC3; mem['h123D]=8'h30; mem['h123E]=8'h12; mem['h123F]=8'hB7;
    mem['h1240]=8'h0E; mem['h1241]=8'hF1; mem['h1242]=8'hF5; mem['h1243]=8'h2A;
    mem['h1244]=8'h9F; mem['h1245]=8'h80; mem['h1246]=8'hEB; mem['h1247]=8'h2A;
    mem['h1248]=8'h08; mem['h1249]=8'h81; mem['h124A]=8'h2F; mem['h124B]=8'h4F;
    mem['h124C]=8'h06; mem['h124D]=8'hFF; mem['h124E]=8'h09; mem['h124F]=8'h23;
    mem['h1250]=8'hCD; mem['h1251]=8'h50; mem['h1252]=8'h07; mem['h1253]=8'hDA;
    mem['h1254]=8'h5D; mem['h1255]=8'h12; mem['h1256]=8'h22; mem['h1257]=8'h08;
    mem['h1258]=8'h81; mem['h1259]=8'h23; mem['h125A]=8'hEB; mem['h125B]=8'hF1;
    mem['h125C]=8'hC9; mem['h125D]=8'hF1; mem['h125E]=8'h1E; mem['h125F]=8'h1A;
    mem['h1260]=8'hCA; mem['h1261]=8'h9C; mem['h1262]=8'h04; mem['h1263]=8'hBF;
    mem['h1264]=8'hF5; mem['h1265]=8'h01; mem['h1266]=8'h41; mem['h1267]=8'h12;
    mem['h1268]=8'hC5; mem['h1269]=8'h2A; mem['h126A]=8'hF4; mem['h126B]=8'h80;
    mem['h126C]=8'h22; mem['h126D]=8'h08; mem['h126E]=8'h81; mem['h126F]=8'h21;
    mem['h1270]=8'h00; mem['h1271]=8'h00; mem['h1272]=8'hE5; mem['h1273]=8'h2A;
    mem['h1274]=8'h9F; mem['h1275]=8'h80; mem['h1276]=8'hE5; mem['h1277]=8'h21;
    mem['h1278]=8'hF8; mem['h1279]=8'h80; mem['h127A]=8'hEB; mem['h127B]=8'h2A;
    mem['h127C]=8'hF6; mem['h127D]=8'h80; mem['h127E]=8'hEB; mem['h127F]=8'hCD;
    mem['h1280]=8'h50; mem['h1281]=8'h07; mem['h1282]=8'h01; mem['h1283]=8'h7A;
    mem['h1284]=8'h12; mem['h1285]=8'hC2; mem['h1286]=8'hCE; mem['h1287]=8'h12;
    mem['h1288]=8'h2A; mem['h1289]=8'h1B; mem['h128A]=8'h81; mem['h128B]=8'hEB;
    mem['h128C]=8'h2A; mem['h128D]=8'h1D; mem['h128E]=8'h81; mem['h128F]=8'hEB;
    mem['h1290]=8'hCD; mem['h1291]=8'h50; mem['h1292]=8'h07; mem['h1293]=8'hCA;
    mem['h1294]=8'hA1; mem['h1295]=8'h12; mem['h1296]=8'h7E; mem['h1297]=8'h23;
    mem['h1298]=8'h23; mem['h1299]=8'hB7; mem['h129A]=8'hCD; mem['h129B]=8'hD1;
    mem['h129C]=8'h12; mem['h129D]=8'hC3; mem['h129E]=8'h8B; mem['h129F]=8'h12;
    mem['h12A0]=8'hC1; mem['h12A1]=8'hEB; mem['h12A2]=8'h2A; mem['h12A3]=8'h1F;
    mem['h12A4]=8'h81; mem['h12A5]=8'hEB; mem['h12A6]=8'hCD; mem['h12A7]=8'h50;
    mem['h12A8]=8'h07; mem['h12A9]=8'hCA; mem['h12AA]=8'hF7; mem['h12AB]=8'h12;
    mem['h12AC]=8'hCD; mem['h12AD]=8'h7E; mem['h12AE]=8'h17; mem['h12AF]=8'h7B;
    mem['h12B0]=8'hE5; mem['h12B1]=8'h09; mem['h12B2]=8'hB7; mem['h12B3]=8'hF2;
    mem['h12B4]=8'hA0; mem['h12B5]=8'h12; mem['h12B6]=8'h22; mem['h12B7]=8'h0A;
    mem['h12B8]=8'h81; mem['h12B9]=8'hE1; mem['h12BA]=8'h4E; mem['h12BB]=8'h06;
    mem['h12BC]=8'h00; mem['h12BD]=8'h09; mem['h12BE]=8'h09; mem['h12BF]=8'h23;
    mem['h12C0]=8'hEB; mem['h12C1]=8'h2A; mem['h12C2]=8'h0A; mem['h12C3]=8'h81;
    mem['h12C4]=8'hEB; mem['h12C5]=8'hCD; mem['h12C6]=8'h50; mem['h12C7]=8'h07;
    mem['h12C8]=8'hCA; mem['h12C9]=8'hA1; mem['h12CA]=8'h12; mem['h12CB]=8'h01;
    mem['h12CC]=8'hC0; mem['h12CD]=8'h12; mem['h12CE]=8'hC5; mem['h12CF]=8'hF6;
    mem['h12D0]=8'h80; mem['h12D1]=8'h7E; mem['h12D2]=8'h23; mem['h12D3]=8'h23;
    mem['h12D4]=8'h5E; mem['h12D5]=8'h23; mem['h12D6]=8'h56; mem['h12D7]=8'h23;
    mem['h12D8]=8'hF0; mem['h12D9]=8'hB7; mem['h12DA]=8'hC8; mem['h12DB]=8'h44;
    mem['h12DC]=8'h4D; mem['h12DD]=8'h2A; mem['h12DE]=8'h08; mem['h12DF]=8'h81;
    mem['h12E0]=8'hCD; mem['h12E1]=8'h50; mem['h12E2]=8'h07; mem['h12E3]=8'h60;
    mem['h12E4]=8'h69; mem['h12E5]=8'hD8; mem['h12E6]=8'hE1; mem['h12E7]=8'hE3;
    mem['h12E8]=8'hCD; mem['h12E9]=8'h50; mem['h12EA]=8'h07; mem['h12EB]=8'hE3;
    mem['h12EC]=8'hE5; mem['h12ED]=8'h60; mem['h12EE]=8'h69; mem['h12EF]=8'hD0;
    mem['h12F0]=8'hC1; mem['h12F1]=8'hF1; mem['h12F2]=8'hF1; mem['h12F3]=8'hE5;
    mem['h12F4]=8'hD5; mem['h12F5]=8'hC5; mem['h12F6]=8'hC9; mem['h12F7]=8'hD1;
    mem['h12F8]=8'hE1; mem['h12F9]=8'h7D; mem['h12FA]=8'hB4; mem['h12FB]=8'hC8;
    mem['h12FC]=8'h2B; mem['h12FD]=8'h46; mem['h12FE]=8'h2B; mem['h12FF]=8'h4E;
    mem['h1300]=8'hE5; mem['h1301]=8'h2B; mem['h1302]=8'h2B; mem['h1303]=8'h6E;
    mem['h1304]=8'h26; mem['h1305]=8'h00; mem['h1306]=8'h09; mem['h1307]=8'h50;
    mem['h1308]=8'h59; mem['h1309]=8'h2B; mem['h130A]=8'h44; mem['h130B]=8'h4D;
    mem['h130C]=8'h2A; mem['h130D]=8'h08; mem['h130E]=8'h81; mem['h130F]=8'hCD;
    mem['h1310]=8'h57; mem['h1311]=8'h04; mem['h1312]=8'hE1; mem['h1313]=8'h71;
    mem['h1314]=8'h23; mem['h1315]=8'h70; mem['h1316]=8'h69; mem['h1317]=8'h60;
    mem['h1318]=8'h2B; mem['h1319]=8'hC3; mem['h131A]=8'h6C; mem['h131B]=8'h12;
    mem['h131C]=8'hC5; mem['h131D]=8'hE5; mem['h131E]=8'h2A; mem['h131F]=8'h29;
    mem['h1320]=8'h81; mem['h1321]=8'hE3; mem['h1322]=8'hCD; mem['h1323]=8'hD6;
    mem['h1324]=8'h0D; mem['h1325]=8'hE3; mem['h1326]=8'hCD; mem['h1327]=8'h51;
    mem['h1328]=8'h0D; mem['h1329]=8'h7E; mem['h132A]=8'hE5; mem['h132B]=8'h2A;
    mem['h132C]=8'h29; mem['h132D]=8'h81; mem['h132E]=8'hE5; mem['h132F]=8'h86;
    mem['h1330]=8'h1E; mem['h1331]=8'h1C; mem['h1332]=8'hDA; mem['h1333]=8'h9C;
    mem['h1334]=8'h04; mem['h1335]=8'hCD; mem['h1336]=8'hD5; mem['h1337]=8'h11;
    mem['h1338]=8'hD1; mem['h1339]=8'hCD; mem['h133A]=8'h6D; mem['h133B]=8'h13;
    mem['h133C]=8'hE3; mem['h133D]=8'hCD; mem['h133E]=8'h6C; mem['h133F]=8'h13;
    mem['h1340]=8'hE5; mem['h1341]=8'h2A; mem['h1342]=8'h06; mem['h1343]=8'h81;
    mem['h1344]=8'hEB; mem['h1345]=8'hCD; mem['h1346]=8'h53; mem['h1347]=8'h13;
    mem['h1348]=8'hCD; mem['h1349]=8'h53; mem['h134A]=8'h13; mem['h134B]=8'h21;
    mem['h134C]=8'h6B; mem['h134D]=8'h0D; mem['h134E]=8'hE3; mem['h134F]=8'hE5;
    mem['h1350]=8'hC3; mem['h1351]=8'h06; mem['h1352]=8'h12; mem['h1353]=8'hE1;
    mem['h1354]=8'hE3; mem['h1355]=8'h7E; mem['h1356]=8'h23; mem['h1357]=8'h23;
    mem['h1358]=8'h4E; mem['h1359]=8'h23; mem['h135A]=8'h46; mem['h135B]=8'h6F;
    mem['h135C]=8'h2C; mem['h135D]=8'h2D; mem['h135E]=8'hC8; mem['h135F]=8'h0A;
    mem['h1360]=8'h12; mem['h1361]=8'h03; mem['h1362]=8'h13; mem['h1363]=8'hC3;
    mem['h1364]=8'h5D; mem['h1365]=8'h13; mem['h1366]=8'hCD; mem['h1367]=8'h51;
    mem['h1368]=8'h0D; mem['h1369]=8'h2A; mem['h136A]=8'h29; mem['h136B]=8'h81;
    mem['h136C]=8'hEB; mem['h136D]=8'hCD; mem['h136E]=8'h87; mem['h136F]=8'h13;
    mem['h1370]=8'hEB; mem['h1371]=8'hC0; mem['h1372]=8'hD5; mem['h1373]=8'h50;
    mem['h1374]=8'h59; mem['h1375]=8'h1B; mem['h1376]=8'h4E; mem['h1377]=8'h2A;
    mem['h1378]=8'h08; mem['h1379]=8'h81; mem['h137A]=8'hCD; mem['h137B]=8'h50;
    mem['h137C]=8'h07; mem['h137D]=8'hC2; mem['h137E]=8'h85; mem['h137F]=8'h13;
    mem['h1380]=8'h47; mem['h1381]=8'h09; mem['h1382]=8'h22; mem['h1383]=8'h08;
    mem['h1384]=8'h81; mem['h1385]=8'hE1; mem['h1386]=8'hC9; mem['h1387]=8'h2A;
    mem['h1388]=8'hF6; mem['h1389]=8'h80; mem['h138A]=8'h2B; mem['h138B]=8'h46;
    mem['h138C]=8'h2B; mem['h138D]=8'h4E; mem['h138E]=8'h2B; mem['h138F]=8'h2B;
    mem['h1390]=8'hCD; mem['h1391]=8'h50; mem['h1392]=8'h07; mem['h1393]=8'hC0;
    mem['h1394]=8'h22; mem['h1395]=8'hF6; mem['h1396]=8'h80; mem['h1397]=8'hC9;
    mem['h1398]=8'h01; mem['h1399]=8'h17; mem['h139A]=8'h11; mem['h139B]=8'hC5;
    mem['h139C]=8'hCD; mem['h139D]=8'h66; mem['h139E]=8'h13; mem['h139F]=8'hAF;
    mem['h13A0]=8'h57; mem['h13A1]=8'h32; mem['h13A2]=8'hF2; mem['h13A3]=8'h80;
    mem['h13A4]=8'h7E; mem['h13A5]=8'hB7; mem['h13A6]=8'hC9; mem['h13A7]=8'h01;
    mem['h13A8]=8'h17; mem['h13A9]=8'h11; mem['h13AA]=8'hC5; mem['h13AB]=8'hCD;
    mem['h13AC]=8'h9C; mem['h13AD]=8'h13; mem['h13AE]=8'hCA; mem['h13AF]=8'hA7;
    mem['h13B0]=8'h09; mem['h13B1]=8'h23; mem['h13B2]=8'h23; mem['h13B3]=8'h5E;
    mem['h13B4]=8'h23; mem['h13B5]=8'h56; mem['h13B6]=8'h1A; mem['h13B7]=8'hC9;
    mem['h13B8]=8'h3E; mem['h13B9]=8'h01; mem['h13BA]=8'hCD; mem['h13BB]=8'hD5;
    mem['h13BC]=8'h11; mem['h13BD]=8'hCD; mem['h13BE]=8'hB1; mem['h13BF]=8'h14;
    mem['h13C0]=8'h2A; mem['h13C1]=8'h06; mem['h13C2]=8'h81; mem['h13C3]=8'h73;
    mem['h13C4]=8'hC1; mem['h13C5]=8'hC3; mem['h13C6]=8'h06; mem['h13C7]=8'h12;
    mem['h13C8]=8'hCD; mem['h13C9]=8'h61; mem['h13CA]=8'h14; mem['h13CB]=8'hAF;
    mem['h13CC]=8'hE3; mem['h13CD]=8'h4F; mem['h13CE]=8'hE5; mem['h13CF]=8'h7E;
    mem['h13D0]=8'hB8; mem['h13D1]=8'hDA; mem['h13D2]=8'hD6; mem['h13D3]=8'h13;
    mem['h13D4]=8'h78; mem['h13D5]=8'h11; mem['h13D6]=8'h0E; mem['h13D7]=8'h00;
    mem['h13D8]=8'hC5; mem['h13D9]=8'hCD; mem['h13DA]=8'h3F; mem['h13DB]=8'h12;
    mem['h13DC]=8'hC1; mem['h13DD]=8'hE1; mem['h13DE]=8'hE5; mem['h13DF]=8'h23;
    mem['h13E0]=8'h23; mem['h13E1]=8'h46; mem['h13E2]=8'h23; mem['h13E3]=8'h66;
    mem['h13E4]=8'h68; mem['h13E5]=8'h06; mem['h13E6]=8'h00; mem['h13E7]=8'h09;
    mem['h13E8]=8'h44; mem['h13E9]=8'h4D; mem['h13EA]=8'hCD; mem['h13EB]=8'hD8;
    mem['h13EC]=8'h11; mem['h13ED]=8'h6F; mem['h13EE]=8'hCD; mem['h13EF]=8'h5C;
    mem['h13F0]=8'h13; mem['h13F1]=8'hD1; mem['h13F2]=8'hCD; mem['h13F3]=8'h6D;
    mem['h13F4]=8'h13; mem['h13F5]=8'hC3; mem['h13F6]=8'h06; mem['h13F7]=8'h12;
    mem['h13F8]=8'hCD; mem['h13F9]=8'h61; mem['h13FA]=8'h14; mem['h13FB]=8'hD1;
    mem['h13FC]=8'hD5; mem['h13FD]=8'h1A; mem['h13FE]=8'h90; mem['h13FF]=8'hC3;
    mem['h1400]=8'hCC; mem['h1401]=8'h13; mem['h1402]=8'hEB; mem['h1403]=8'h7E;
    mem['h1404]=8'hCD; mem['h1405]=8'h66; mem['h1406]=8'h14; mem['h1407]=8'h04;
    mem['h1408]=8'h05; mem['h1409]=8'hCA; mem['h140A]=8'hA7; mem['h140B]=8'h09;
    mem['h140C]=8'hC5; mem['h140D]=8'h1E; mem['h140E]=8'hFF; mem['h140F]=8'hFE;
    mem['h1410]=8'h29; mem['h1411]=8'hCA; mem['h1412]=8'h1B; mem['h1413]=8'h14;
    mem['h1414]=8'hCD; mem['h1415]=8'h56; mem['h1416]=8'h07; mem['h1417]=8'h2C;
    mem['h1418]=8'hCD; mem['h1419]=8'hAE; mem['h141A]=8'h14; mem['h141B]=8'hCD;
    mem['h141C]=8'h56; mem['h141D]=8'h07; mem['h141E]=8'h29; mem['h141F]=8'hF1;
    mem['h1420]=8'hE3; mem['h1421]=8'h01; mem['h1422]=8'hCE; mem['h1423]=8'h13;
    mem['h1424]=8'hC5; mem['h1425]=8'h3D; mem['h1426]=8'hBE; mem['h1427]=8'h06;
    mem['h1428]=8'h00; mem['h1429]=8'hD0; mem['h142A]=8'h4F; mem['h142B]=8'h7E;
    mem['h142C]=8'h91; mem['h142D]=8'hBB; mem['h142E]=8'h47; mem['h142F]=8'hD8;
    mem['h1430]=8'h43; mem['h1431]=8'hC9; mem['h1432]=8'hCD; mem['h1433]=8'h9C;
    mem['h1434]=8'h13; mem['h1435]=8'hCA; mem['h1436]=8'h4F; mem['h1437]=8'h15;
    mem['h1438]=8'h5F; mem['h1439]=8'h23; mem['h143A]=8'h23; mem['h143B]=8'h7E;
    mem['h143C]=8'h23; mem['h143D]=8'h66; mem['h143E]=8'h6F; mem['h143F]=8'hE5;
    mem['h1440]=8'h19; mem['h1441]=8'h46; mem['h1442]=8'h72; mem['h1443]=8'hE3;
    mem['h1444]=8'hC5; mem['h1445]=8'h7E; mem['h1446]=8'hFE; mem['h1447]=8'h24;
    mem['h1448]=8'hC2; mem['h1449]=8'h50; mem['h144A]=8'h14; mem['h144B]=8'hCD;
    mem['h144C]=8'h7A; mem['h144D]=8'h1C; mem['h144E]=8'h18; mem['h144F]=8'h0D;
    mem['h1450]=8'hFE; mem['h1451]=8'h25; mem['h1452]=8'hC2; mem['h1453]=8'h5A;
    mem['h1454]=8'h14; mem['h1455]=8'hCD; mem['h1456]=8'hEA; mem['h1457]=8'h1C;
    mem['h1458]=8'h18; mem['h1459]=8'h03; mem['h145A]=8'hCD; mem['h145B]=8'h36;
    mem['h145C]=8'h18; mem['h145D]=8'hC1; mem['h145E]=8'hE1; mem['h145F]=8'h70;
    mem['h1460]=8'hC9; mem['h1461]=8'hEB; mem['h1462]=8'hCD; mem['h1463]=8'h56;
    mem['h1464]=8'h07; mem['h1465]=8'h29; mem['h1466]=8'hC1; mem['h1467]=8'hD1;
    mem['h1468]=8'hC5; mem['h1469]=8'h43; mem['h146A]=8'hC9; mem['h146B]=8'hCD;
    mem['h146C]=8'hB1; mem['h146D]=8'h14; mem['h146E]=8'h32; mem['h146F]=8'h84;
    mem['h1470]=8'h80; mem['h1471]=8'hCD; mem['h1472]=8'h83; mem['h1473]=8'h80;
    mem['h1474]=8'hC3; mem['h1475]=8'h17; mem['h1476]=8'h11; mem['h1477]=8'hCD;
    mem['h1478]=8'h9B; mem['h1479]=8'h14; mem['h147A]=8'hC3; mem['h147B]=8'h4B;
    mem['h147C]=8'h80; mem['h147D]=8'hCD; mem['h147E]=8'h9B; mem['h147F]=8'h14;
    mem['h1480]=8'hF5; mem['h1481]=8'h1E; mem['h1482]=8'h00; mem['h1483]=8'h2B;
    mem['h1484]=8'hCD; mem['h1485]=8'hE0; mem['h1486]=8'h08; mem['h1487]=8'hCA;
    mem['h1488]=8'h91; mem['h1489]=8'h14; mem['h148A]=8'hCD; mem['h148B]=8'h56;
    mem['h148C]=8'h07; mem['h148D]=8'h2C; mem['h148E]=8'hCD; mem['h148F]=8'hAE;
    mem['h1490]=8'h14; mem['h1491]=8'hC1; mem['h1492]=8'hCD; mem['h1493]=8'h83;
    mem['h1494]=8'h80; mem['h1495]=8'hAB; mem['h1496]=8'hA0; mem['h1497]=8'hCA;
    mem['h1498]=8'h92; mem['h1499]=8'h14; mem['h149A]=8'hC9; mem['h149B]=8'hCD;
    mem['h149C]=8'hAE; mem['h149D]=8'h14; mem['h149E]=8'h32; mem['h149F]=8'h84;
    mem['h14A0]=8'h80; mem['h14A1]=8'h32; mem['h14A2]=8'h4C; mem['h14A3]=8'h80;
    mem['h14A4]=8'hCD; mem['h14A5]=8'h56; mem['h14A6]=8'h07; mem['h14A7]=8'h2C;
    mem['h14A8]=8'hC3; mem['h14A9]=8'hAE; mem['h14AA]=8'h14; mem['h14AB]=8'hCD;
    mem['h14AC]=8'hE0; mem['h14AD]=8'h08; mem['h14AE]=8'hCD; mem['h14AF]=8'h4D;
    mem['h14B0]=8'h0D; mem['h14B1]=8'hCD; mem['h14B2]=8'h8C; mem['h14B3]=8'h09;
    mem['h14B4]=8'h7A; mem['h14B5]=8'hB7; mem['h14B6]=8'hC2; mem['h14B7]=8'hA7;
    mem['h14B8]=8'h09; mem['h14B9]=8'h2B; mem['h14BA]=8'hCD; mem['h14BB]=8'hE0;
    mem['h14BC]=8'h08; mem['h14BD]=8'h7B; mem['h14BE]=8'hC9; mem['h14BF]=8'hCD;
    mem['h14C0]=8'h92; mem['h14C1]=8'h09; mem['h14C2]=8'h1A; mem['h14C3]=8'hC3;
    mem['h14C4]=8'h17; mem['h14C5]=8'h11; mem['h14C6]=8'hCD; mem['h14C7]=8'h4D;
    mem['h14C8]=8'h0D; mem['h14C9]=8'hCD; mem['h14CA]=8'h92; mem['h14CB]=8'h09;
    mem['h14CC]=8'hD5; mem['h14CD]=8'hCD; mem['h14CE]=8'h56; mem['h14CF]=8'h07;
    mem['h14D0]=8'h2C; mem['h14D1]=8'hCD; mem['h14D2]=8'hAE; mem['h14D3]=8'h14;
    mem['h14D4]=8'hD1; mem['h14D5]=8'h12; mem['h14D6]=8'hC9; mem['h14D7]=8'h21;
    mem['h14D8]=8'hAD; mem['h14D9]=8'h19; mem['h14DA]=8'hCD; mem['h14DB]=8'h7E;
    mem['h14DC]=8'h17; mem['h14DD]=8'hC3; mem['h14DE]=8'hE9; mem['h14DF]=8'h14;
    mem['h14E0]=8'hCD; mem['h14E1]=8'h7E; mem['h14E2]=8'h17; mem['h14E3]=8'h21;
    mem['h14E4]=8'hC1; mem['h14E5]=8'hD1; mem['h14E6]=8'hCD; mem['h14E7]=8'h58;
    mem['h14E8]=8'h17; mem['h14E9]=8'h78; mem['h14EA]=8'hB7; mem['h14EB]=8'hC8;
    mem['h14EC]=8'h3A; mem['h14ED]=8'h2C; mem['h14EE]=8'h81; mem['h14EF]=8'hB7;
    mem['h14F0]=8'hCA; mem['h14F1]=8'h70; mem['h14F2]=8'h17; mem['h14F3]=8'h90;
    mem['h14F4]=8'hD2; mem['h14F5]=8'h03; mem['h14F6]=8'h15; mem['h14F7]=8'h2F;
    mem['h14F8]=8'h3C; mem['h14F9]=8'hEB; mem['h14FA]=8'hCD; mem['h14FB]=8'h60;
    mem['h14FC]=8'h17; mem['h14FD]=8'hEB; mem['h14FE]=8'hCD; mem['h14FF]=8'h70;
    mem['h1500]=8'h17; mem['h1501]=8'hC1; mem['h1502]=8'hD1; mem['h1503]=8'hFE;
    mem['h1504]=8'h19; mem['h1505]=8'hD0; mem['h1506]=8'hF5; mem['h1507]=8'hCD;
    mem['h1508]=8'h95; mem['h1509]=8'h17; mem['h150A]=8'h67; mem['h150B]=8'hF1;
    mem['h150C]=8'hCD; mem['h150D]=8'hAE; mem['h150E]=8'h15; mem['h150F]=8'hB4;
    mem['h1510]=8'h21; mem['h1511]=8'h29; mem['h1512]=8'h81; mem['h1513]=8'hF2;
    mem['h1514]=8'h29; mem['h1515]=8'h15; mem['h1516]=8'hCD; mem['h1517]=8'h8E;
    mem['h1518]=8'h15; mem['h1519]=8'hD2; mem['h151A]=8'h6F; mem['h151B]=8'h15;
    mem['h151C]=8'h23; mem['h151D]=8'h34; mem['h151E]=8'hCA; mem['h151F]=8'h97;
    mem['h1520]=8'h04; mem['h1521]=8'h2E; mem['h1522]=8'h01; mem['h1523]=8'hCD;
    mem['h1524]=8'hC4; mem['h1525]=8'h15; mem['h1526]=8'hC3; mem['h1527]=8'h6F;
    mem['h1528]=8'h15; mem['h1529]=8'hAF; mem['h152A]=8'h90; mem['h152B]=8'h47;
    mem['h152C]=8'h7E; mem['h152D]=8'h9B; mem['h152E]=8'h5F; mem['h152F]=8'h23;
    mem['h1530]=8'h7E; mem['h1531]=8'h9A; mem['h1532]=8'h57; mem['h1533]=8'h23;
    mem['h1534]=8'h7E; mem['h1535]=8'h99; mem['h1536]=8'h4F; mem['h1537]=8'hDC;
    mem['h1538]=8'h9A; mem['h1539]=8'h15; mem['h153A]=8'h68; mem['h153B]=8'h63;
    mem['h153C]=8'hAF; mem['h153D]=8'h47; mem['h153E]=8'h79; mem['h153F]=8'hB7;
    mem['h1540]=8'hC2; mem['h1541]=8'h5C; mem['h1542]=8'h15; mem['h1543]=8'h4A;
    mem['h1544]=8'h54; mem['h1545]=8'h65; mem['h1546]=8'h6F; mem['h1547]=8'h78;
    mem['h1548]=8'hD6; mem['h1549]=8'h08; mem['h154A]=8'hFE; mem['h154B]=8'hE0;
    mem['h154C]=8'hC2; mem['h154D]=8'h3D; mem['h154E]=8'h15; mem['h154F]=8'hAF;
    mem['h1550]=8'h32; mem['h1551]=8'h2C; mem['h1552]=8'h81; mem['h1553]=8'hC9;
    mem['h1554]=8'h05; mem['h1555]=8'h29; mem['h1556]=8'h7A; mem['h1557]=8'h17;
    mem['h1558]=8'h57; mem['h1559]=8'h79; mem['h155A]=8'h8F; mem['h155B]=8'h4F;
    mem['h155C]=8'hF2; mem['h155D]=8'h54; mem['h155E]=8'h15; mem['h155F]=8'h78;
    mem['h1560]=8'h5C; mem['h1561]=8'h45; mem['h1562]=8'hB7; mem['h1563]=8'hCA;
    mem['h1564]=8'h6F; mem['h1565]=8'h15; mem['h1566]=8'h21; mem['h1567]=8'h2C;
    mem['h1568]=8'h81; mem['h1569]=8'h86; mem['h156A]=8'h77; mem['h156B]=8'hD2;
    mem['h156C]=8'h4F; mem['h156D]=8'h15; mem['h156E]=8'hC8; mem['h156F]=8'h78;
    mem['h1570]=8'h21; mem['h1571]=8'h2C; mem['h1572]=8'h81; mem['h1573]=8'hB7;
    mem['h1574]=8'hFC; mem['h1575]=8'h81; mem['h1576]=8'h15; mem['h1577]=8'h46;
    mem['h1578]=8'h23; mem['h1579]=8'h7E; mem['h157A]=8'hE6; mem['h157B]=8'h80;
    mem['h157C]=8'hA9; mem['h157D]=8'h4F; mem['h157E]=8'hC3; mem['h157F]=8'h70;
    mem['h1580]=8'h17; mem['h1581]=8'h1C; mem['h1582]=8'hC0; mem['h1583]=8'h14;
    mem['h1584]=8'hC0; mem['h1585]=8'h0C; mem['h1586]=8'hC0; mem['h1587]=8'h0E;
    mem['h1588]=8'h80; mem['h1589]=8'h34; mem['h158A]=8'hC0; mem['h158B]=8'hC3;
    mem['h158C]=8'h97; mem['h158D]=8'h04; mem['h158E]=8'h7E; mem['h158F]=8'h83;
    mem['h1590]=8'h5F; mem['h1591]=8'h23; mem['h1592]=8'h7E; mem['h1593]=8'h8A;
    mem['h1594]=8'h57; mem['h1595]=8'h23; mem['h1596]=8'h7E; mem['h1597]=8'h89;
    mem['h1598]=8'h4F; mem['h1599]=8'hC9; mem['h159A]=8'h21; mem['h159B]=8'h2D;
    mem['h159C]=8'h81; mem['h159D]=8'h7E; mem['h159E]=8'h2F; mem['h159F]=8'h77;
    mem['h15A0]=8'hAF; mem['h15A1]=8'h6F; mem['h15A2]=8'h90; mem['h15A3]=8'h47;
    mem['h15A4]=8'h7D; mem['h15A5]=8'h9B; mem['h15A6]=8'h5F; mem['h15A7]=8'h7D;
    mem['h15A8]=8'h9A; mem['h15A9]=8'h57; mem['h15AA]=8'h7D; mem['h15AB]=8'h99;
    mem['h15AC]=8'h4F; mem['h15AD]=8'hC9; mem['h15AE]=8'h06; mem['h15AF]=8'h00;
    mem['h15B0]=8'hD6; mem['h15B1]=8'h08; mem['h15B2]=8'hDA; mem['h15B3]=8'hBD;
    mem['h15B4]=8'h15; mem['h15B5]=8'h43; mem['h15B6]=8'h5A; mem['h15B7]=8'h51;
    mem['h15B8]=8'h0E; mem['h15B9]=8'h00; mem['h15BA]=8'hC3; mem['h15BB]=8'hB0;
    mem['h15BC]=8'h15; mem['h15BD]=8'hC6; mem['h15BE]=8'h09; mem['h15BF]=8'h6F;
    mem['h15C0]=8'hAF; mem['h15C1]=8'h2D; mem['h15C2]=8'hC8; mem['h15C3]=8'h79;
    mem['h15C4]=8'h1F; mem['h15C5]=8'h4F; mem['h15C6]=8'h7A; mem['h15C7]=8'h1F;
    mem['h15C8]=8'h57; mem['h15C9]=8'h7B; mem['h15CA]=8'h1F; mem['h15CB]=8'h5F;
    mem['h15CC]=8'h78; mem['h15CD]=8'h1F; mem['h15CE]=8'h47; mem['h15CF]=8'hC3;
    mem['h15D0]=8'hC0; mem['h15D1]=8'h15; mem['h15D2]=8'h00; mem['h15D3]=8'h00;
    mem['h15D4]=8'h00; mem['h15D5]=8'h81; mem['h15D6]=8'h03; mem['h15D7]=8'hAA;
    mem['h15D8]=8'h56; mem['h15D9]=8'h19; mem['h15DA]=8'h80; mem['h15DB]=8'hF1;
    mem['h15DC]=8'h22; mem['h15DD]=8'h76; mem['h15DE]=8'h80; mem['h15DF]=8'h45;
    mem['h15E0]=8'hAA; mem['h15E1]=8'h38; mem['h15E2]=8'h82; mem['h15E3]=8'hCD;
    mem['h15E4]=8'h2F; mem['h15E5]=8'h17; mem['h15E6]=8'hB7; mem['h15E7]=8'hEA;
    mem['h15E8]=8'hA7; mem['h15E9]=8'h09; mem['h15EA]=8'h21; mem['h15EB]=8'h2C;
    mem['h15EC]=8'h81; mem['h15ED]=8'h7E; mem['h15EE]=8'h01; mem['h15EF]=8'h35;
    mem['h15F0]=8'h80; mem['h15F1]=8'h11; mem['h15F2]=8'hF3; mem['h15F3]=8'h04;
    mem['h15F4]=8'h90; mem['h15F5]=8'hF5; mem['h15F6]=8'h70; mem['h15F7]=8'hD5;
    mem['h15F8]=8'hC5; mem['h15F9]=8'hCD; mem['h15FA]=8'hE9; mem['h15FB]=8'h14;
    mem['h15FC]=8'hC1; mem['h15FD]=8'hD1; mem['h15FE]=8'h04; mem['h15FF]=8'hCD;
    mem['h1600]=8'h85; mem['h1601]=8'h16; mem['h1602]=8'h21; mem['h1603]=8'hD2;
    mem['h1604]=8'h15; mem['h1605]=8'hCD; mem['h1606]=8'hE0; mem['h1607]=8'h14;
    mem['h1608]=8'h21; mem['h1609]=8'hD6; mem['h160A]=8'h15; mem['h160B]=8'hCD;
    mem['h160C]=8'h77; mem['h160D]=8'h1A; mem['h160E]=8'h01; mem['h160F]=8'h80;
    mem['h1610]=8'h80; mem['h1611]=8'h11; mem['h1612]=8'h00; mem['h1613]=8'h00;
    mem['h1614]=8'hCD; mem['h1615]=8'hE9; mem['h1616]=8'h14; mem['h1617]=8'hF1;
    mem['h1618]=8'hCD; mem['h1619]=8'hAA; mem['h161A]=8'h18; mem['h161B]=8'h01;
    mem['h161C]=8'h31; mem['h161D]=8'h80; mem['h161E]=8'h11; mem['h161F]=8'h18;
    mem['h1620]=8'h72; mem['h1621]=8'h21; mem['h1622]=8'hC1; mem['h1623]=8'hD1;
    mem['h1624]=8'hCD; mem['h1625]=8'h2F; mem['h1626]=8'h17; mem['h1627]=8'hC8;
    mem['h1628]=8'h2E; mem['h1629]=8'h00; mem['h162A]=8'hCD; mem['h162B]=8'hED;
    mem['h162C]=8'h16; mem['h162D]=8'h79; mem['h162E]=8'h32; mem['h162F]=8'h3B;
    mem['h1630]=8'h81; mem['h1631]=8'hEB; mem['h1632]=8'h22; mem['h1633]=8'h3C;
    mem['h1634]=8'h81; mem['h1635]=8'h01; mem['h1636]=8'h00; mem['h1637]=8'h00;
    mem['h1638]=8'h50; mem['h1639]=8'h58; mem['h163A]=8'h21; mem['h163B]=8'h3A;
    mem['h163C]=8'h15; mem['h163D]=8'hE5; mem['h163E]=8'h21; mem['h163F]=8'h46;
    mem['h1640]=8'h16; mem['h1641]=8'hE5; mem['h1642]=8'hE5; mem['h1643]=8'h21;
    mem['h1644]=8'h29; mem['h1645]=8'h81; mem['h1646]=8'h7E; mem['h1647]=8'h23;
    mem['h1648]=8'hB7; mem['h1649]=8'hCA; mem['h164A]=8'h72; mem['h164B]=8'h16;
    mem['h164C]=8'hE5; mem['h164D]=8'h2E; mem['h164E]=8'h08; mem['h164F]=8'h1F;
    mem['h1650]=8'h67; mem['h1651]=8'h79; mem['h1652]=8'hD2; mem['h1653]=8'h60;
    mem['h1654]=8'h16; mem['h1655]=8'hE5; mem['h1656]=8'h2A; mem['h1657]=8'h3C;
    mem['h1658]=8'h81; mem['h1659]=8'h19; mem['h165A]=8'hEB; mem['h165B]=8'hE1;
    mem['h165C]=8'h3A; mem['h165D]=8'h3B; mem['h165E]=8'h81; mem['h165F]=8'h89;
    mem['h1660]=8'h1F; mem['h1661]=8'h4F; mem['h1662]=8'h7A; mem['h1663]=8'h1F;
    mem['h1664]=8'h57; mem['h1665]=8'h7B; mem['h1666]=8'h1F; mem['h1667]=8'h5F;
    mem['h1668]=8'h78; mem['h1669]=8'h1F; mem['h166A]=8'h47; mem['h166B]=8'h2D;
    mem['h166C]=8'h7C; mem['h166D]=8'hC2; mem['h166E]=8'h4F; mem['h166F]=8'h16;
    mem['h1670]=8'hE1; mem['h1671]=8'hC9; mem['h1672]=8'h43; mem['h1673]=8'h5A;
    mem['h1674]=8'h51; mem['h1675]=8'h4F; mem['h1676]=8'hC9; mem['h1677]=8'hCD;
    mem['h1678]=8'h60; mem['h1679]=8'h17; mem['h167A]=8'h01; mem['h167B]=8'h20;
    mem['h167C]=8'h84; mem['h167D]=8'h11; mem['h167E]=8'h00; mem['h167F]=8'h00;
    mem['h1680]=8'hCD; mem['h1681]=8'h70; mem['h1682]=8'h17; mem['h1683]=8'hC1;
    mem['h1684]=8'hD1; mem['h1685]=8'hCD; mem['h1686]=8'h2F; mem['h1687]=8'h17;
    mem['h1688]=8'hCA; mem['h1689]=8'h8B; mem['h168A]=8'h04; mem['h168B]=8'h2E;
    mem['h168C]=8'hFF; mem['h168D]=8'hCD; mem['h168E]=8'hED; mem['h168F]=8'h16;
    mem['h1690]=8'h34; mem['h1691]=8'h34; mem['h1692]=8'h2B; mem['h1693]=8'h7E;
    mem['h1694]=8'h32; mem['h1695]=8'h57; mem['h1696]=8'h80; mem['h1697]=8'h2B;
    mem['h1698]=8'h7E; mem['h1699]=8'h32; mem['h169A]=8'h53; mem['h169B]=8'h80;
    mem['h169C]=8'h2B; mem['h169D]=8'h7E; mem['h169E]=8'h32; mem['h169F]=8'h4F;
    mem['h16A0]=8'h80; mem['h16A1]=8'h41; mem['h16A2]=8'hEB; mem['h16A3]=8'hAF;
    mem['h16A4]=8'h4F; mem['h16A5]=8'h57; mem['h16A6]=8'h5F; mem['h16A7]=8'h32;
    mem['h16A8]=8'h5A; mem['h16A9]=8'h80; mem['h16AA]=8'hE5; mem['h16AB]=8'hC5;
    mem['h16AC]=8'h7D; mem['h16AD]=8'hCD; mem['h16AE]=8'h4E; mem['h16AF]=8'h80;
    mem['h16B0]=8'hDE; mem['h16B1]=8'h00; mem['h16B2]=8'h3F; mem['h16B3]=8'hD2;
    mem['h16B4]=8'hBD; mem['h16B5]=8'h16; mem['h16B6]=8'h32; mem['h16B7]=8'h5A;
    mem['h16B8]=8'h80; mem['h16B9]=8'hF1; mem['h16BA]=8'hF1; mem['h16BB]=8'h37;
    mem['h16BC]=8'hD2; mem['h16BD]=8'hC1; mem['h16BE]=8'hE1; mem['h16BF]=8'h79;
    mem['h16C0]=8'h3C; mem['h16C1]=8'h3D; mem['h16C2]=8'h1F; mem['h16C3]=8'hFA;
    mem['h16C4]=8'h70; mem['h16C5]=8'h15; mem['h16C6]=8'h17; mem['h16C7]=8'h7B;
    mem['h16C8]=8'h17; mem['h16C9]=8'h5F; mem['h16CA]=8'h7A; mem['h16CB]=8'h17;
    mem['h16CC]=8'h57; mem['h16CD]=8'h79; mem['h16CE]=8'h17; mem['h16CF]=8'h4F;
    mem['h16D0]=8'h29; mem['h16D1]=8'h78; mem['h16D2]=8'h17; mem['h16D3]=8'h47;
    mem['h16D4]=8'h3A; mem['h16D5]=8'h5A; mem['h16D6]=8'h80; mem['h16D7]=8'h17;
    mem['h16D8]=8'h32; mem['h16D9]=8'h5A; mem['h16DA]=8'h80; mem['h16DB]=8'h79;
    mem['h16DC]=8'hB2; mem['h16DD]=8'hB3; mem['h16DE]=8'hC2; mem['h16DF]=8'hAA;
    mem['h16E0]=8'h16; mem['h16E1]=8'hE5; mem['h16E2]=8'h21; mem['h16E3]=8'h2C;
    mem['h16E4]=8'h81; mem['h16E5]=8'h35; mem['h16E6]=8'hE1; mem['h16E7]=8'hC2;
    mem['h16E8]=8'hAA; mem['h16E9]=8'h16; mem['h16EA]=8'hC3; mem['h16EB]=8'h97;
    mem['h16EC]=8'h04; mem['h16ED]=8'h78; mem['h16EE]=8'hB7; mem['h16EF]=8'hCA;
    mem['h16F0]=8'h11; mem['h16F1]=8'h17; mem['h16F2]=8'h7D; mem['h16F3]=8'h21;
    mem['h16F4]=8'h2C; mem['h16F5]=8'h81; mem['h16F6]=8'hAE; mem['h16F7]=8'h80;
    mem['h16F8]=8'h47; mem['h16F9]=8'h1F; mem['h16FA]=8'hA8; mem['h16FB]=8'h78;
    mem['h16FC]=8'hF2; mem['h16FD]=8'h10; mem['h16FE]=8'h17; mem['h16FF]=8'hC6;
    mem['h1700]=8'h80; mem['h1701]=8'h77; mem['h1702]=8'hCA; mem['h1703]=8'h70;
    mem['h1704]=8'h16; mem['h1705]=8'hCD; mem['h1706]=8'h95; mem['h1707]=8'h17;
    mem['h1708]=8'h77; mem['h1709]=8'h2B; mem['h170A]=8'hC9; mem['h170B]=8'hCD;
    mem['h170C]=8'h2F; mem['h170D]=8'h17; mem['h170E]=8'h2F; mem['h170F]=8'hE1;
    mem['h1710]=8'hB7; mem['h1711]=8'hE1; mem['h1712]=8'hF2; mem['h1713]=8'h4F;
    mem['h1714]=8'h15; mem['h1715]=8'hC3; mem['h1716]=8'h97; mem['h1717]=8'h04;
    mem['h1718]=8'hCD; mem['h1719]=8'h7B; mem['h171A]=8'h17; mem['h171B]=8'h78;
    mem['h171C]=8'hB7; mem['h171D]=8'hC8; mem['h171E]=8'hC6; mem['h171F]=8'h02;
    mem['h1720]=8'hDA; mem['h1721]=8'h97; mem['h1722]=8'h04; mem['h1723]=8'h47;
    mem['h1724]=8'hCD; mem['h1725]=8'hE9; mem['h1726]=8'h14; mem['h1727]=8'h21;
    mem['h1728]=8'h2C; mem['h1729]=8'h81; mem['h172A]=8'h34; mem['h172B]=8'hC0;
    mem['h172C]=8'hC3; mem['h172D]=8'h97; mem['h172E]=8'h04; mem['h172F]=8'h3A;
    mem['h1730]=8'h2C; mem['h1731]=8'h81; mem['h1732]=8'hB7; mem['h1733]=8'hC8;
    mem['h1734]=8'h3A; mem['h1735]=8'h2B; mem['h1736]=8'h81; mem['h1737]=8'hFE;
    mem['h1738]=8'h2F; mem['h1739]=8'h17; mem['h173A]=8'h9F; mem['h173B]=8'hC0;
    mem['h173C]=8'h3C; mem['h173D]=8'hC9; mem['h173E]=8'hCD; mem['h173F]=8'h2F;
    mem['h1740]=8'h17; mem['h1741]=8'h06; mem['h1742]=8'h88; mem['h1743]=8'h11;
    mem['h1744]=8'h00; mem['h1745]=8'h00; mem['h1746]=8'h21; mem['h1747]=8'h2C;
    mem['h1748]=8'h81; mem['h1749]=8'h4F; mem['h174A]=8'h70; mem['h174B]=8'h06;
    mem['h174C]=8'h00; mem['h174D]=8'h23; mem['h174E]=8'h36; mem['h174F]=8'h80;
    mem['h1750]=8'h17; mem['h1751]=8'hC3; mem['h1752]=8'h37; mem['h1753]=8'h15;
    mem['h1754]=8'hCD; mem['h1755]=8'h2F; mem['h1756]=8'h17; mem['h1757]=8'hF0;
    mem['h1758]=8'h21; mem['h1759]=8'h2B; mem['h175A]=8'h81; mem['h175B]=8'h7E;
    mem['h175C]=8'hEE; mem['h175D]=8'h80; mem['h175E]=8'h77; mem['h175F]=8'hC9;
    mem['h1760]=8'hEB; mem['h1761]=8'h2A; mem['h1762]=8'h29; mem['h1763]=8'h81;
    mem['h1764]=8'hE3; mem['h1765]=8'hE5; mem['h1766]=8'h2A; mem['h1767]=8'h2B;
    mem['h1768]=8'h81; mem['h1769]=8'hE3; mem['h176A]=8'hE5; mem['h176B]=8'hEB;
    mem['h176C]=8'hC9; mem['h176D]=8'hCD; mem['h176E]=8'h7E; mem['h176F]=8'h17;
    mem['h1770]=8'hEB; mem['h1771]=8'h22; mem['h1772]=8'h29; mem['h1773]=8'h81;
    mem['h1774]=8'h60; mem['h1775]=8'h69; mem['h1776]=8'h22; mem['h1777]=8'h2B;
    mem['h1778]=8'h81; mem['h1779]=8'hEB; mem['h177A]=8'hC9; mem['h177B]=8'h21;
    mem['h177C]=8'h29; mem['h177D]=8'h81; mem['h177E]=8'h5E; mem['h177F]=8'h23;
    mem['h1780]=8'h56; mem['h1781]=8'h23; mem['h1782]=8'h4E; mem['h1783]=8'h23;
    mem['h1784]=8'h46; mem['h1785]=8'h23; mem['h1786]=8'hC9; mem['h1787]=8'h11;
    mem['h1788]=8'h29; mem['h1789]=8'h81; mem['h178A]=8'h06; mem['h178B]=8'h04;
    mem['h178C]=8'h1A; mem['h178D]=8'h77; mem['h178E]=8'h13; mem['h178F]=8'h23;
    mem['h1790]=8'h05; mem['h1791]=8'hC2; mem['h1792]=8'h8C; mem['h1793]=8'h17;
    mem['h1794]=8'hC9; mem['h1795]=8'h21; mem['h1796]=8'h2B; mem['h1797]=8'h81;
    mem['h1798]=8'h7E; mem['h1799]=8'h07; mem['h179A]=8'h37; mem['h179B]=8'h1F;
    mem['h179C]=8'h77; mem['h179D]=8'h3F; mem['h179E]=8'h1F; mem['h179F]=8'h23;
    mem['h17A0]=8'h23; mem['h17A1]=8'h77; mem['h17A2]=8'h79; mem['h17A3]=8'h07;
    mem['h17A4]=8'h37; mem['h17A5]=8'h1F; mem['h17A6]=8'h4F; mem['h17A7]=8'h1F;
    mem['h17A8]=8'hAE; mem['h17A9]=8'hC9; mem['h17AA]=8'h78; mem['h17AB]=8'hB7;
    mem['h17AC]=8'hCA; mem['h17AD]=8'h2F; mem['h17AE]=8'h17; mem['h17AF]=8'h21;
    mem['h17B0]=8'h38; mem['h17B1]=8'h17; mem['h17B2]=8'hE5; mem['h17B3]=8'hCD;
    mem['h17B4]=8'h2F; mem['h17B5]=8'h17; mem['h17B6]=8'h79; mem['h17B7]=8'hC8;
    mem['h17B8]=8'h21; mem['h17B9]=8'h2B; mem['h17BA]=8'h81; mem['h17BB]=8'hAE;
    mem['h17BC]=8'h79; mem['h17BD]=8'hF8; mem['h17BE]=8'hCD; mem['h17BF]=8'hC4;
    mem['h17C0]=8'h17; mem['h17C1]=8'h1F; mem['h17C2]=8'hA9; mem['h17C3]=8'hC9;
    mem['h17C4]=8'h23; mem['h17C5]=8'h78; mem['h17C6]=8'hBE; mem['h17C7]=8'hC0;
    mem['h17C8]=8'h2B; mem['h17C9]=8'h79; mem['h17CA]=8'hBE; mem['h17CB]=8'hC0;
    mem['h17CC]=8'h2B; mem['h17CD]=8'h7A; mem['h17CE]=8'hBE; mem['h17CF]=8'hC0;
    mem['h17D0]=8'h2B; mem['h17D1]=8'h7B; mem['h17D2]=8'h96; mem['h17D3]=8'hC0;
    mem['h17D4]=8'hE1; mem['h17D5]=8'hE1; mem['h17D6]=8'hC9; mem['h17D7]=8'h47;
    mem['h17D8]=8'h4F; mem['h17D9]=8'h57; mem['h17DA]=8'h5F; mem['h17DB]=8'hB7;
    mem['h17DC]=8'hC8; mem['h17DD]=8'hE5; mem['h17DE]=8'hCD; mem['h17DF]=8'h7B;
    mem['h17E0]=8'h17; mem['h17E1]=8'hCD; mem['h17E2]=8'h95; mem['h17E3]=8'h17;
    mem['h17E4]=8'hAE; mem['h17E5]=8'h67; mem['h17E6]=8'hFC; mem['h17E7]=8'hFB;
    mem['h17E8]=8'h17; mem['h17E9]=8'h3E; mem['h17EA]=8'h98; mem['h17EB]=8'h90;
    mem['h17EC]=8'hCD; mem['h17ED]=8'hAE; mem['h17EE]=8'h15; mem['h17EF]=8'h7C;
    mem['h17F0]=8'h17; mem['h17F1]=8'hDC; mem['h17F2]=8'h81; mem['h17F3]=8'h15;
    mem['h17F4]=8'h06; mem['h17F5]=8'h00; mem['h17F6]=8'hDC; mem['h17F7]=8'h9A;
    mem['h17F8]=8'h15; mem['h17F9]=8'hE1; mem['h17FA]=8'hC9; mem['h17FB]=8'h1B;
    mem['h17FC]=8'h7A; mem['h17FD]=8'hA3; mem['h17FE]=8'h3C; mem['h17FF]=8'hC0;
    mem['h1800]=8'h0B; mem['h1801]=8'hC9; mem['h1802]=8'h21; mem['h1803]=8'h2C;
    mem['h1804]=8'h81; mem['h1805]=8'h7E; mem['h1806]=8'hFE; mem['h1807]=8'h98;
    mem['h1808]=8'h3A; mem['h1809]=8'h29; mem['h180A]=8'h81; mem['h180B]=8'hD0;
    mem['h180C]=8'h7E; mem['h180D]=8'hCD; mem['h180E]=8'hD7; mem['h180F]=8'h17;
    mem['h1810]=8'h36; mem['h1811]=8'h98; mem['h1812]=8'h7B; mem['h1813]=8'hF5;
    mem['h1814]=8'h79; mem['h1815]=8'h17; mem['h1816]=8'hCD; mem['h1817]=8'h37;
    mem['h1818]=8'h15; mem['h1819]=8'hF1; mem['h181A]=8'hC9; mem['h181B]=8'h21;
    mem['h181C]=8'h00; mem['h181D]=8'h00; mem['h181E]=8'h78; mem['h181F]=8'hB1;
    mem['h1820]=8'hC8; mem['h1821]=8'h3E; mem['h1822]=8'h10; mem['h1823]=8'h29;
    mem['h1824]=8'hDA; mem['h1825]=8'h5B; mem['h1826]=8'h10; mem['h1827]=8'hEB;
    mem['h1828]=8'h29; mem['h1829]=8'hEB; mem['h182A]=8'hD2; mem['h182B]=8'h31;
    mem['h182C]=8'h18; mem['h182D]=8'h09; mem['h182E]=8'hDA; mem['h182F]=8'h5B;
    mem['h1830]=8'h10; mem['h1831]=8'h3D; mem['h1832]=8'hC2; mem['h1833]=8'h23;
    mem['h1834]=8'h18; mem['h1835]=8'hC9; mem['h1836]=8'hFE; mem['h1837]=8'h2D;
    mem['h1838]=8'hF5; mem['h1839]=8'hCA; mem['h183A]=8'h42; mem['h183B]=8'h18;
    mem['h183C]=8'hFE; mem['h183D]=8'h2B; mem['h183E]=8'hCA; mem['h183F]=8'h42;
    mem['h1840]=8'h18; mem['h1841]=8'h2B; mem['h1842]=8'hCD; mem['h1843]=8'h4F;
    mem['h1844]=8'h15; mem['h1845]=8'h47; mem['h1846]=8'h57; mem['h1847]=8'h5F;
    mem['h1848]=8'h2F; mem['h1849]=8'h4F; mem['h184A]=8'hCD; mem['h184B]=8'hE0;
    mem['h184C]=8'h08; mem['h184D]=8'hDA; mem['h184E]=8'h93; mem['h184F]=8'h18;
    mem['h1850]=8'hFE; mem['h1851]=8'h2E; mem['h1852]=8'hCA; mem['h1853]=8'h6E;
    mem['h1854]=8'h18; mem['h1855]=8'hFE; mem['h1856]=8'h45; mem['h1857]=8'hC2;
    mem['h1858]=8'h72; mem['h1859]=8'h18; mem['h185A]=8'hCD; mem['h185B]=8'hE0;
    mem['h185C]=8'h08; mem['h185D]=8'hCD; mem['h185E]=8'h86; mem['h185F]=8'h0E;
    mem['h1860]=8'hCD; mem['h1861]=8'hE0; mem['h1862]=8'h08; mem['h1863]=8'hDA;
    mem['h1864]=8'hB5; mem['h1865]=8'h18; mem['h1866]=8'h14; mem['h1867]=8'hC2;
    mem['h1868]=8'h72; mem['h1869]=8'h18; mem['h186A]=8'hAF; mem['h186B]=8'h93;
    mem['h186C]=8'h5F; mem['h186D]=8'h0C; mem['h186E]=8'h0C; mem['h186F]=8'hCA;
    mem['h1870]=8'h4A; mem['h1871]=8'h18; mem['h1872]=8'hE5; mem['h1873]=8'h7B;
    mem['h1874]=8'h90; mem['h1875]=8'hF4; mem['h1876]=8'h8B; mem['h1877]=8'h18;
    mem['h1878]=8'hF2; mem['h1879]=8'h81; mem['h187A]=8'h18; mem['h187B]=8'hF5;
    mem['h187C]=8'hCD; mem['h187D]=8'h77; mem['h187E]=8'h16; mem['h187F]=8'hF1;
    mem['h1880]=8'h3C; mem['h1881]=8'hC2; mem['h1882]=8'h75; mem['h1883]=8'h18;
    mem['h1884]=8'hD1; mem['h1885]=8'hF1; mem['h1886]=8'hCC; mem['h1887]=8'h58;
    mem['h1888]=8'h17; mem['h1889]=8'hEB; mem['h188A]=8'hC9; mem['h188B]=8'hC8;
    mem['h188C]=8'hF5; mem['h188D]=8'hCD; mem['h188E]=8'h18; mem['h188F]=8'h17;
    mem['h1890]=8'hF1; mem['h1891]=8'h3D; mem['h1892]=8'hC9; mem['h1893]=8'hD5;
    mem['h1894]=8'h57; mem['h1895]=8'h78; mem['h1896]=8'h89; mem['h1897]=8'h47;
    mem['h1898]=8'hC5; mem['h1899]=8'hE5; mem['h189A]=8'hD5; mem['h189B]=8'hCD;
    mem['h189C]=8'h18; mem['h189D]=8'h17; mem['h189E]=8'hF1; mem['h189F]=8'hD6;
    mem['h18A0]=8'h30; mem['h18A1]=8'hCD; mem['h18A2]=8'hAA; mem['h18A3]=8'h18;
    mem['h18A4]=8'hE1; mem['h18A5]=8'hC1; mem['h18A6]=8'hD1; mem['h18A7]=8'hC3;
    mem['h18A8]=8'h4A; mem['h18A9]=8'h18; mem['h18AA]=8'hCD; mem['h18AB]=8'h60;
    mem['h18AC]=8'h17; mem['h18AD]=8'hCD; mem['h18AE]=8'h41; mem['h18AF]=8'h17;
    mem['h18B0]=8'hC1; mem['h18B1]=8'hD1; mem['h18B2]=8'hC3; mem['h18B3]=8'hE9;
    mem['h18B4]=8'h14; mem['h18B5]=8'h7B; mem['h18B6]=8'h07; mem['h18B7]=8'h07;
    mem['h18B8]=8'h83; mem['h18B9]=8'h07; mem['h18BA]=8'h86; mem['h18BB]=8'hD6;
    mem['h18BC]=8'h30; mem['h18BD]=8'h5F; mem['h18BE]=8'hC3; mem['h18BF]=8'h60;
    mem['h18C0]=8'h18; mem['h18C1]=8'hE5; mem['h18C2]=8'h21; mem['h18C3]=8'h20;
    mem['h18C4]=8'h04; mem['h18C5]=8'hCD; mem['h18C6]=8'h26; mem['h18C7]=8'h12;
    mem['h18C8]=8'hE1; mem['h18C9]=8'hEB; mem['h18CA]=8'hAF; mem['h18CB]=8'h06;
    mem['h18CC]=8'h98; mem['h18CD]=8'hCD; mem['h18CE]=8'h46; mem['h18CF]=8'h17;
    mem['h18D0]=8'h21; mem['h18D1]=8'h25; mem['h18D2]=8'h12; mem['h18D3]=8'hE5;
    mem['h18D4]=8'h21; mem['h18D5]=8'h2E; mem['h18D6]=8'h81; mem['h18D7]=8'hE5;
    mem['h18D8]=8'hCD; mem['h18D9]=8'h2F; mem['h18DA]=8'h17; mem['h18DB]=8'h36;
    mem['h18DC]=8'h20; mem['h18DD]=8'hF2; mem['h18DE]=8'hE2; mem['h18DF]=8'h18;
    mem['h18E0]=8'h36; mem['h18E1]=8'h2D; mem['h18E2]=8'h23; mem['h18E3]=8'h36;
    mem['h18E4]=8'h30; mem['h18E5]=8'hCA; mem['h18E6]=8'h98; mem['h18E7]=8'h19;
    mem['h18E8]=8'hE5; mem['h18E9]=8'hFC; mem['h18EA]=8'h58; mem['h18EB]=8'h17;
    mem['h18EC]=8'hAF; mem['h18ED]=8'hF5; mem['h18EE]=8'hCD; mem['h18EF]=8'h9E;
    mem['h18F0]=8'h19; mem['h18F1]=8'h01; mem['h18F2]=8'h43; mem['h18F3]=8'h91;
    mem['h18F4]=8'h11; mem['h18F5]=8'hF8; mem['h18F6]=8'h4F; mem['h18F7]=8'hCD;
    mem['h18F8]=8'hAA; mem['h18F9]=8'h17; mem['h18FA]=8'hB7; mem['h18FB]=8'hE2;
    mem['h18FC]=8'h0F; mem['h18FD]=8'h19; mem['h18FE]=8'hF1; mem['h18FF]=8'hCD;
    mem['h1900]=8'h8C; mem['h1901]=8'h18; mem['h1902]=8'hF5; mem['h1903]=8'hC3;
    mem['h1904]=8'hF1; mem['h1905]=8'h18; mem['h1906]=8'hCD; mem['h1907]=8'h77;
    mem['h1908]=8'h16; mem['h1909]=8'hF1; mem['h190A]=8'h3C; mem['h190B]=8'hF5;
    mem['h190C]=8'hCD; mem['h190D]=8'h9E; mem['h190E]=8'h19; mem['h190F]=8'hCD;
    mem['h1910]=8'hD7; mem['h1911]=8'h14; mem['h1912]=8'h3C; mem['h1913]=8'hCD;
    mem['h1914]=8'hD7; mem['h1915]=8'h17; mem['h1916]=8'hCD; mem['h1917]=8'h70;
    mem['h1918]=8'h17; mem['h1919]=8'h01; mem['h191A]=8'h06; mem['h191B]=8'h03;
    mem['h191C]=8'hF1; mem['h191D]=8'h81; mem['h191E]=8'h3C; mem['h191F]=8'hFA;
    mem['h1920]=8'h2B; mem['h1921]=8'h19; mem['h1922]=8'hFE; mem['h1923]=8'h08;
    mem['h1924]=8'hD2; mem['h1925]=8'h2B; mem['h1926]=8'h19; mem['h1927]=8'h3C;
    mem['h1928]=8'h47; mem['h1929]=8'h3E; mem['h192A]=8'h02; mem['h192B]=8'h3D;
    mem['h192C]=8'h3D; mem['h192D]=8'hE1; mem['h192E]=8'hF5; mem['h192F]=8'h11;
    mem['h1930]=8'hB1; mem['h1931]=8'h19; mem['h1932]=8'h05; mem['h1933]=8'hC2;
    mem['h1934]=8'h3C; mem['h1935]=8'h19; mem['h1936]=8'h36; mem['h1937]=8'h2E;
    mem['h1938]=8'h23; mem['h1939]=8'h36; mem['h193A]=8'h30; mem['h193B]=8'h23;
    mem['h193C]=8'h05; mem['h193D]=8'h36; mem['h193E]=8'h2E; mem['h193F]=8'hCC;
    mem['h1940]=8'h85; mem['h1941]=8'h17; mem['h1942]=8'hC5; mem['h1943]=8'hE5;
    mem['h1944]=8'hD5; mem['h1945]=8'hCD; mem['h1946]=8'h7B; mem['h1947]=8'h17;
    mem['h1948]=8'hE1; mem['h1949]=8'h06; mem['h194A]=8'h2F; mem['h194B]=8'h04;
    mem['h194C]=8'h7B; mem['h194D]=8'h96; mem['h194E]=8'h5F; mem['h194F]=8'h23;
    mem['h1950]=8'h7A; mem['h1951]=8'h9E; mem['h1952]=8'h57; mem['h1953]=8'h23;
    mem['h1954]=8'h79; mem['h1955]=8'h9E; mem['h1956]=8'h4F; mem['h1957]=8'h2B;
    mem['h1958]=8'h2B; mem['h1959]=8'hD2; mem['h195A]=8'h4B; mem['h195B]=8'h19;
    mem['h195C]=8'hCD; mem['h195D]=8'h8E; mem['h195E]=8'h15; mem['h195F]=8'h23;
    mem['h1960]=8'hCD; mem['h1961]=8'h70; mem['h1962]=8'h17; mem['h1963]=8'hEB;
    mem['h1964]=8'hE1; mem['h1965]=8'h70; mem['h1966]=8'h23; mem['h1967]=8'hC1;
    mem['h1968]=8'h0D; mem['h1969]=8'hC2; mem['h196A]=8'h3C; mem['h196B]=8'h19;
    mem['h196C]=8'h05; mem['h196D]=8'hCA; mem['h196E]=8'h7C; mem['h196F]=8'h19;
    mem['h1970]=8'h2B; mem['h1971]=8'h7E; mem['h1972]=8'hFE; mem['h1973]=8'h30;
    mem['h1974]=8'hCA; mem['h1975]=8'h70; mem['h1976]=8'h19; mem['h1977]=8'hFE;
    mem['h1978]=8'h2E; mem['h1979]=8'hC4; mem['h197A]=8'h85; mem['h197B]=8'h17;
    mem['h197C]=8'hF1; mem['h197D]=8'hCA; mem['h197E]=8'h9B; mem['h197F]=8'h19;
    mem['h1980]=8'h36; mem['h1981]=8'h45; mem['h1982]=8'h23; mem['h1983]=8'h36;
    mem['h1984]=8'h2B; mem['h1985]=8'hF2; mem['h1986]=8'h8C; mem['h1987]=8'h19;
    mem['h1988]=8'h36; mem['h1989]=8'h2D; mem['h198A]=8'h2F; mem['h198B]=8'h3C;
    mem['h198C]=8'h06; mem['h198D]=8'h2F; mem['h198E]=8'h04; mem['h198F]=8'hD6;
    mem['h1990]=8'h0A; mem['h1991]=8'hD2; mem['h1992]=8'h8E; mem['h1993]=8'h19;
    mem['h1994]=8'hC6; mem['h1995]=8'h3A; mem['h1996]=8'h23; mem['h1997]=8'h70;
    mem['h1998]=8'h23; mem['h1999]=8'h77; mem['h199A]=8'h23; mem['h199B]=8'h71;
    mem['h199C]=8'hE1; mem['h199D]=8'hC9; mem['h199E]=8'h01; mem['h199F]=8'h74;
    mem['h19A0]=8'h94; mem['h19A1]=8'h11; mem['h19A2]=8'hF7; mem['h19A3]=8'h23;
    mem['h19A4]=8'hCD; mem['h19A5]=8'hAA; mem['h19A6]=8'h17; mem['h19A7]=8'hB7;
    mem['h19A8]=8'hE1; mem['h19A9]=8'hE2; mem['h19AA]=8'h06; mem['h19AB]=8'h19;
    mem['h19AC]=8'hE9; mem['h19AD]=8'h00; mem['h19AE]=8'h00; mem['h19AF]=8'h00;
    mem['h19B0]=8'h80; mem['h19B1]=8'hA0; mem['h19B2]=8'h86; mem['h19B3]=8'h01;
    mem['h19B4]=8'h10; mem['h19B5]=8'h27; mem['h19B6]=8'h00; mem['h19B7]=8'hE8;
    mem['h19B8]=8'h03; mem['h19B9]=8'h00; mem['h19BA]=8'h64; mem['h19BB]=8'h00;
    mem['h19BC]=8'h00; mem['h19BD]=8'h0A; mem['h19BE]=8'h00; mem['h19BF]=8'h00;
    mem['h19C0]=8'h01; mem['h19C1]=8'h00; mem['h19C2]=8'h00; mem['h19C3]=8'h21;
    mem['h19C4]=8'h58; mem['h19C5]=8'h17; mem['h19C6]=8'hE3; mem['h19C7]=8'hE9;
    mem['h19C8]=8'hCD; mem['h19C9]=8'h60; mem['h19CA]=8'h17; mem['h19CB]=8'h21;
    mem['h19CC]=8'hAD; mem['h19CD]=8'h19; mem['h19CE]=8'hCD; mem['h19CF]=8'h6D;
    mem['h19D0]=8'h17; mem['h19D1]=8'hC1; mem['h19D2]=8'hD1; mem['h19D3]=8'hCD;
    mem['h19D4]=8'h2F; mem['h19D5]=8'h17; mem['h19D6]=8'h78; mem['h19D7]=8'hCA;
    mem['h19D8]=8'h16; mem['h19D9]=8'h1A; mem['h19DA]=8'hF2; mem['h19DB]=8'hE1;
    mem['h19DC]=8'h19; mem['h19DD]=8'hB7; mem['h19DE]=8'hCA; mem['h19DF]=8'h8B;
    mem['h19E0]=8'h04; mem['h19E1]=8'hB7; mem['h19E2]=8'hCA; mem['h19E3]=8'h50;
    mem['h19E4]=8'h15; mem['h19E5]=8'hD5; mem['h19E6]=8'hC5; mem['h19E7]=8'h79;
    mem['h19E8]=8'hF6; mem['h19E9]=8'h7F; mem['h19EA]=8'hCD; mem['h19EB]=8'h7B;
    mem['h19EC]=8'h17; mem['h19ED]=8'hF2; mem['h19EE]=8'hFE; mem['h19EF]=8'h19;
    mem['h19F0]=8'hD5; mem['h19F1]=8'hC5; mem['h19F2]=8'hCD; mem['h19F3]=8'h02;
    mem['h19F4]=8'h18; mem['h19F5]=8'hC1; mem['h19F6]=8'hD1; mem['h19F7]=8'hF5;
    mem['h19F8]=8'hCD; mem['h19F9]=8'hAA; mem['h19FA]=8'h17; mem['h19FB]=8'hE1;
    mem['h19FC]=8'h7C; mem['h19FD]=8'h1F; mem['h19FE]=8'hE1; mem['h19FF]=8'h22;
    mem['h1A00]=8'h2B; mem['h1A01]=8'h81; mem['h1A02]=8'hE1; mem['h1A03]=8'h22;
    mem['h1A04]=8'h29; mem['h1A05]=8'h81; mem['h1A06]=8'hDC; mem['h1A07]=8'hC3;
    mem['h1A08]=8'h19; mem['h1A09]=8'hCC; mem['h1A0A]=8'h58; mem['h1A0B]=8'h17;
    mem['h1A0C]=8'hD5; mem['h1A0D]=8'hC5; mem['h1A0E]=8'hCD; mem['h1A0F]=8'hE3;
    mem['h1A10]=8'h15; mem['h1A11]=8'hC1; mem['h1A12]=8'hD1; mem['h1A13]=8'hCD;
    mem['h1A14]=8'h24; mem['h1A15]=8'h16; mem['h1A16]=8'hCD; mem['h1A17]=8'h60;
    mem['h1A18]=8'h17; mem['h1A19]=8'h01; mem['h1A1A]=8'h38; mem['h1A1B]=8'h81;
    mem['h1A1C]=8'h11; mem['h1A1D]=8'h3B; mem['h1A1E]=8'hAA; mem['h1A1F]=8'hCD;
    mem['h1A20]=8'h24; mem['h1A21]=8'h16; mem['h1A22]=8'h3A; mem['h1A23]=8'h2C;
    mem['h1A24]=8'h81; mem['h1A25]=8'hFE; mem['h1A26]=8'h88; mem['h1A27]=8'hD2;
    mem['h1A28]=8'h0B; mem['h1A29]=8'h17; mem['h1A2A]=8'hCD; mem['h1A2B]=8'h02;
    mem['h1A2C]=8'h18; mem['h1A2D]=8'hC6; mem['h1A2E]=8'h80; mem['h1A2F]=8'hC6;
    mem['h1A30]=8'h02; mem['h1A31]=8'hDA; mem['h1A32]=8'h0B; mem['h1A33]=8'h17;
    mem['h1A34]=8'hF5; mem['h1A35]=8'h21; mem['h1A36]=8'hD2; mem['h1A37]=8'h15;
    mem['h1A38]=8'hCD; mem['h1A39]=8'hDA; mem['h1A3A]=8'h14; mem['h1A3B]=8'hCD;
    mem['h1A3C]=8'h1B; mem['h1A3D]=8'h16; mem['h1A3E]=8'hF1; mem['h1A3F]=8'hC1;
    mem['h1A40]=8'hD1; mem['h1A41]=8'hF5; mem['h1A42]=8'hCD; mem['h1A43]=8'hE6;
    mem['h1A44]=8'h14; mem['h1A45]=8'hCD; mem['h1A46]=8'h58; mem['h1A47]=8'h17;
    mem['h1A48]=8'h21; mem['h1A49]=8'h56; mem['h1A4A]=8'h1A; mem['h1A4B]=8'hCD;
    mem['h1A4C]=8'h86; mem['h1A4D]=8'h1A; mem['h1A4E]=8'h11; mem['h1A4F]=8'h00;
    mem['h1A50]=8'h00; mem['h1A51]=8'hC1; mem['h1A52]=8'h4A; mem['h1A53]=8'hC3;
    mem['h1A54]=8'h24; mem['h1A55]=8'h16; mem['h1A56]=8'h08; mem['h1A57]=8'h40;
    mem['h1A58]=8'h2E; mem['h1A59]=8'h94; mem['h1A5A]=8'h74; mem['h1A5B]=8'h70;
    mem['h1A5C]=8'h4F; mem['h1A5D]=8'h2E; mem['h1A5E]=8'h77; mem['h1A5F]=8'h6E;
    mem['h1A60]=8'h02; mem['h1A61]=8'h88; mem['h1A62]=8'h7A; mem['h1A63]=8'hE6;
    mem['h1A64]=8'hA0; mem['h1A65]=8'h2A; mem['h1A66]=8'h7C; mem['h1A67]=8'h50;
    mem['h1A68]=8'hAA; mem['h1A69]=8'hAA; mem['h1A6A]=8'h7E; mem['h1A6B]=8'hFF;
    mem['h1A6C]=8'hFF; mem['h1A6D]=8'h7F; mem['h1A6E]=8'h7F; mem['h1A6F]=8'h00;
    mem['h1A70]=8'h00; mem['h1A71]=8'h80; mem['h1A72]=8'h81; mem['h1A73]=8'h00;
    mem['h1A74]=8'h00; mem['h1A75]=8'h00; mem['h1A76]=8'h81; mem['h1A77]=8'hCD;
    mem['h1A78]=8'h60; mem['h1A79]=8'h17; mem['h1A7A]=8'h11; mem['h1A7B]=8'h22;
    mem['h1A7C]=8'h16; mem['h1A7D]=8'hD5; mem['h1A7E]=8'hE5; mem['h1A7F]=8'hCD;
    mem['h1A80]=8'h7B; mem['h1A81]=8'h17; mem['h1A82]=8'hCD; mem['h1A83]=8'h24;
    mem['h1A84]=8'h16; mem['h1A85]=8'hE1; mem['h1A86]=8'hCD; mem['h1A87]=8'h60;
    mem['h1A88]=8'h17; mem['h1A89]=8'h7E; mem['h1A8A]=8'h23; mem['h1A8B]=8'hCD;
    mem['h1A8C]=8'h6D; mem['h1A8D]=8'h17; mem['h1A8E]=8'h06; mem['h1A8F]=8'hF1;
    mem['h1A90]=8'hC1; mem['h1A91]=8'hD1; mem['h1A92]=8'h3D; mem['h1A93]=8'hC8;
    mem['h1A94]=8'hD5; mem['h1A95]=8'hC5; mem['h1A96]=8'hF5; mem['h1A97]=8'hE5;
    mem['h1A98]=8'hCD; mem['h1A99]=8'h24; mem['h1A9A]=8'h16; mem['h1A9B]=8'hE1;
    mem['h1A9C]=8'hCD; mem['h1A9D]=8'h7E; mem['h1A9E]=8'h17; mem['h1A9F]=8'hE5;
    mem['h1AA0]=8'hCD; mem['h1AA1]=8'hE9; mem['h1AA2]=8'h14; mem['h1AA3]=8'hE1;
    mem['h1AA4]=8'hC3; mem['h1AA5]=8'h8F; mem['h1AA6]=8'h1A; mem['h1AA7]=8'hCD;
    mem['h1AA8]=8'h2F; mem['h1AA9]=8'h17; mem['h1AAA]=8'h21; mem['h1AAB]=8'h5E;
    mem['h1AAC]=8'h80; mem['h1AAD]=8'hFA; mem['h1AAE]=8'h08; mem['h1AAF]=8'h1B;
    mem['h1AB0]=8'h21; mem['h1AB1]=8'h7F; mem['h1AB2]=8'h80; mem['h1AB3]=8'hCD;
    mem['h1AB4]=8'h6D; mem['h1AB5]=8'h17; mem['h1AB6]=8'h21; mem['h1AB7]=8'h5E;
    mem['h1AB8]=8'h80; mem['h1AB9]=8'hC8; mem['h1ABA]=8'h86; mem['h1ABB]=8'hE6;
    mem['h1ABC]=8'h07; mem['h1ABD]=8'h06; mem['h1ABE]=8'h00; mem['h1ABF]=8'h77;
    mem['h1AC0]=8'h23; mem['h1AC1]=8'h87; mem['h1AC2]=8'h87; mem['h1AC3]=8'h4F;
    mem['h1AC4]=8'h09; mem['h1AC5]=8'hCD; mem['h1AC6]=8'h7E; mem['h1AC7]=8'h17;
    mem['h1AC8]=8'hCD; mem['h1AC9]=8'h24; mem['h1ACA]=8'h16; mem['h1ACB]=8'h3A;
    mem['h1ACC]=8'h5D; mem['h1ACD]=8'h80; mem['h1ACE]=8'h3C; mem['h1ACF]=8'hE6;
    mem['h1AD0]=8'h03; mem['h1AD1]=8'h06; mem['h1AD2]=8'h00; mem['h1AD3]=8'hFE;
    mem['h1AD4]=8'h01; mem['h1AD5]=8'h88; mem['h1AD6]=8'h32; mem['h1AD7]=8'h5D;
    mem['h1AD8]=8'h80; mem['h1AD9]=8'h21; mem['h1ADA]=8'h0C; mem['h1ADB]=8'h1B;
    mem['h1ADC]=8'h87; mem['h1ADD]=8'h87; mem['h1ADE]=8'h4F; mem['h1ADF]=8'h09;
    mem['h1AE0]=8'hCD; mem['h1AE1]=8'hDA; mem['h1AE2]=8'h14; mem['h1AE3]=8'hCD;
    mem['h1AE4]=8'h7B; mem['h1AE5]=8'h17; mem['h1AE6]=8'h7B; mem['h1AE7]=8'h59;
    mem['h1AE8]=8'hEE; mem['h1AE9]=8'h4F; mem['h1AEA]=8'h4F; mem['h1AEB]=8'h36;
    mem['h1AEC]=8'h80; mem['h1AED]=8'h2B; mem['h1AEE]=8'h46; mem['h1AEF]=8'h36;
    mem['h1AF0]=8'h80; mem['h1AF1]=8'h21; mem['h1AF2]=8'h5C; mem['h1AF3]=8'h80;
    mem['h1AF4]=8'h34; mem['h1AF5]=8'h7E; mem['h1AF6]=8'hD6; mem['h1AF7]=8'hAB;
    mem['h1AF8]=8'hC2; mem['h1AF9]=8'hFF; mem['h1AFA]=8'h1A; mem['h1AFB]=8'h77;
    mem['h1AFC]=8'h0C; mem['h1AFD]=8'h15; mem['h1AFE]=8'h1C; mem['h1AFF]=8'hCD;
    mem['h1B00]=8'h3A; mem['h1B01]=8'h15; mem['h1B02]=8'h21; mem['h1B03]=8'h7F;
    mem['h1B04]=8'h80; mem['h1B05]=8'hC3; mem['h1B06]=8'h87; mem['h1B07]=8'h17;
    mem['h1B08]=8'h77; mem['h1B09]=8'h2B; mem['h1B0A]=8'h77; mem['h1B0B]=8'h2B;
    mem['h1B0C]=8'h77; mem['h1B0D]=8'hC3; mem['h1B0E]=8'hE3; mem['h1B0F]=8'h1A;
    mem['h1B10]=8'h68; mem['h1B11]=8'hB1; mem['h1B12]=8'h46; mem['h1B13]=8'h68;
    mem['h1B14]=8'h99; mem['h1B15]=8'hE9; mem['h1B16]=8'h92; mem['h1B17]=8'h69;
    mem['h1B18]=8'h10; mem['h1B19]=8'hD1; mem['h1B1A]=8'h75; mem['h1B1B]=8'h68;
    mem['h1B1C]=8'h21; mem['h1B1D]=8'h66; mem['h1B1E]=8'h1B; mem['h1B1F]=8'hCD;
    mem['h1B20]=8'hDA; mem['h1B21]=8'h14; mem['h1B22]=8'hCD; mem['h1B23]=8'h60;
    mem['h1B24]=8'h17; mem['h1B25]=8'h01; mem['h1B26]=8'h49; mem['h1B27]=8'h83;
    mem['h1B28]=8'h11; mem['h1B29]=8'hDB; mem['h1B2A]=8'h0F; mem['h1B2B]=8'hCD;
    mem['h1B2C]=8'h70; mem['h1B2D]=8'h17; mem['h1B2E]=8'hC1; mem['h1B2F]=8'hD1;
    mem['h1B30]=8'hCD; mem['h1B31]=8'h85; mem['h1B32]=8'h16; mem['h1B33]=8'hCD;
    mem['h1B34]=8'h60; mem['h1B35]=8'h17; mem['h1B36]=8'hCD; mem['h1B37]=8'h02;
    mem['h1B38]=8'h18; mem['h1B39]=8'hC1; mem['h1B3A]=8'hD1; mem['h1B3B]=8'hCD;
    mem['h1B3C]=8'hE6; mem['h1B3D]=8'h14; mem['h1B3E]=8'h21; mem['h1B3F]=8'h6A;
    mem['h1B40]=8'h1B; mem['h1B41]=8'hCD; mem['h1B42]=8'hE0; mem['h1B43]=8'h14;
    mem['h1B44]=8'hCD; mem['h1B45]=8'h2F; mem['h1B46]=8'h17; mem['h1B47]=8'h37;
    mem['h1B48]=8'hF2; mem['h1B49]=8'h52; mem['h1B4A]=8'h1B; mem['h1B4B]=8'hCD;
    mem['h1B4C]=8'hD7; mem['h1B4D]=8'h14; mem['h1B4E]=8'hCD; mem['h1B4F]=8'h2F;
    mem['h1B50]=8'h17; mem['h1B51]=8'hB7; mem['h1B52]=8'hF5; mem['h1B53]=8'hF4;
    mem['h1B54]=8'h58; mem['h1B55]=8'h17; mem['h1B56]=8'h21; mem['h1B57]=8'h6A;
    mem['h1B58]=8'h1B; mem['h1B59]=8'hCD; mem['h1B5A]=8'hDA; mem['h1B5B]=8'h14;
    mem['h1B5C]=8'hF1; mem['h1B5D]=8'hD4; mem['h1B5E]=8'h58; mem['h1B5F]=8'h17;
    mem['h1B60]=8'h21; mem['h1B61]=8'h6E; mem['h1B62]=8'h1B; mem['h1B63]=8'hC3;
    mem['h1B64]=8'h77; mem['h1B65]=8'h1A; mem['h1B66]=8'hDB; mem['h1B67]=8'h0F;
    mem['h1B68]=8'h49; mem['h1B69]=8'h81; mem['h1B6A]=8'h00; mem['h1B6B]=8'h00;
    mem['h1B6C]=8'h00; mem['h1B6D]=8'h7F; mem['h1B6E]=8'h05; mem['h1B6F]=8'hBA;
    mem['h1B70]=8'hD7; mem['h1B71]=8'h1E; mem['h1B72]=8'h86; mem['h1B73]=8'h64;
    mem['h1B74]=8'h26; mem['h1B75]=8'h99; mem['h1B76]=8'h87; mem['h1B77]=8'h58;
    mem['h1B78]=8'h34; mem['h1B79]=8'h23; mem['h1B7A]=8'h87; mem['h1B7B]=8'hE0;
    mem['h1B7C]=8'h5D; mem['h1B7D]=8'hA5; mem['h1B7E]=8'h86; mem['h1B7F]=8'hDA;
    mem['h1B80]=8'h0F; mem['h1B81]=8'h49; mem['h1B82]=8'h83; mem['h1B83]=8'hCD;
    mem['h1B84]=8'h60; mem['h1B85]=8'h17; mem['h1B86]=8'hCD; mem['h1B87]=8'h22;
    mem['h1B88]=8'h1B; mem['h1B89]=8'hC1; mem['h1B8A]=8'hE1; mem['h1B8B]=8'hCD;
    mem['h1B8C]=8'h60; mem['h1B8D]=8'h17; mem['h1B8E]=8'hEB; mem['h1B8F]=8'hCD;
    mem['h1B90]=8'h70; mem['h1B91]=8'h17; mem['h1B92]=8'hCD; mem['h1B93]=8'h1C;
    mem['h1B94]=8'h1B; mem['h1B95]=8'hC3; mem['h1B96]=8'h83; mem['h1B97]=8'h16;
    mem['h1B98]=8'hCD; mem['h1B99]=8'h2F; mem['h1B9A]=8'h17; mem['h1B9B]=8'hFC;
    mem['h1B9C]=8'hC3; mem['h1B9D]=8'h19; mem['h1B9E]=8'hFC; mem['h1B9F]=8'h58;
    mem['h1BA0]=8'h17; mem['h1BA1]=8'h3A; mem['h1BA2]=8'h2C; mem['h1BA3]=8'h81;
    mem['h1BA4]=8'hFE; mem['h1BA5]=8'h81; mem['h1BA6]=8'hDA; mem['h1BA7]=8'hB5;
    mem['h1BA8]=8'h1B; mem['h1BA9]=8'h01; mem['h1BAA]=8'h00; mem['h1BAB]=8'h81;
    mem['h1BAC]=8'h51; mem['h1BAD]=8'h59; mem['h1BAE]=8'hCD; mem['h1BAF]=8'h85;
    mem['h1BB0]=8'h16; mem['h1BB1]=8'h21; mem['h1BB2]=8'hE0; mem['h1BB3]=8'h14;
    mem['h1BB4]=8'hE5; mem['h1BB5]=8'h21; mem['h1BB6]=8'hBF; mem['h1BB7]=8'h1B;
    mem['h1BB8]=8'hCD; mem['h1BB9]=8'h77; mem['h1BBA]=8'h1A; mem['h1BBB]=8'h21;
    mem['h1BBC]=8'h66; mem['h1BBD]=8'h1B; mem['h1BBE]=8'hC9; mem['h1BBF]=8'h09;
    mem['h1BC0]=8'h4A; mem['h1BC1]=8'hD7; mem['h1BC2]=8'h3B; mem['h1BC3]=8'h78;
    mem['h1BC4]=8'h02; mem['h1BC5]=8'h6E; mem['h1BC6]=8'h84; mem['h1BC7]=8'h7B;
    mem['h1BC8]=8'hFE; mem['h1BC9]=8'hC1; mem['h1BCA]=8'h2F; mem['h1BCB]=8'h7C;
    mem['h1BCC]=8'h74; mem['h1BCD]=8'h31; mem['h1BCE]=8'h9A; mem['h1BCF]=8'h7D;
    mem['h1BD0]=8'h84; mem['h1BD1]=8'h3D; mem['h1BD2]=8'h5A; mem['h1BD3]=8'h7D;
    mem['h1BD4]=8'hC8; mem['h1BD5]=8'h7F; mem['h1BD6]=8'h91; mem['h1BD7]=8'h7E;
    mem['h1BD8]=8'hE4; mem['h1BD9]=8'hBB; mem['h1BDA]=8'h4C; mem['h1BDB]=8'h7E;
    mem['h1BDC]=8'h6C; mem['h1BDD]=8'hAA; mem['h1BDE]=8'hAA; mem['h1BDF]=8'h7F;
    mem['h1BE0]=8'h00; mem['h1BE1]=8'h00; mem['h1BE2]=8'h00; mem['h1BE3]=8'h81;
    mem['h1BE4]=8'hC9; mem['h1BE5]=8'hD7; mem['h1BE6]=8'hC9; mem['h1BE7]=8'h3E;
    mem['h1BE8]=8'h0C; mem['h1BE9]=8'hC3; mem['h1BEA]=8'h1D; mem['h1BEB]=8'h1D;
    mem['h1BEC]=8'hCD; mem['h1BED]=8'hAE; mem['h1BEE]=8'h14; mem['h1BEF]=8'h7B;
    mem['h1BF0]=8'h32; mem['h1BF1]=8'h87; mem['h1BF2]=8'h80; mem['h1BF3]=8'hC9;
    mem['h1BF4]=8'hCD; mem['h1BF5]=8'h4D; mem['h1BF6]=8'h0D; mem['h1BF7]=8'hCD;
    mem['h1BF8]=8'h92; mem['h1BF9]=8'h09; mem['h1BFA]=8'hED; mem['h1BFB]=8'h53;
    mem['h1BFC]=8'h8B; mem['h1BFD]=8'h80; mem['h1BFE]=8'hED; mem['h1BFF]=8'h53;
    mem['h1C00]=8'h8D; mem['h1C01]=8'h80; mem['h1C02]=8'hC9; mem['h1C03]=8'hCD;
    mem['h1C04]=8'h92; mem['h1C05]=8'h09; mem['h1C06]=8'hD5; mem['h1C07]=8'hE1;
    mem['h1C08]=8'h46; mem['h1C09]=8'h23; mem['h1C0A]=8'h7E; mem['h1C0B]=8'hC3;
    mem['h1C0C]=8'h08; mem['h1C0D]=8'h11; mem['h1C0E]=8'hCD; mem['h1C0F]=8'h4D;
    mem['h1C10]=8'h0D; mem['h1C11]=8'hCD; mem['h1C12]=8'h92; mem['h1C13]=8'h09;
    mem['h1C14]=8'hD5; mem['h1C15]=8'hCD; mem['h1C16]=8'h56; mem['h1C17]=8'h07;
    mem['h1C18]=8'h2C; mem['h1C19]=8'hCD; mem['h1C1A]=8'h4D; mem['h1C1B]=8'h0D;
    mem['h1C1C]=8'hCD; mem['h1C1D]=8'h92; mem['h1C1E]=8'h09; mem['h1C1F]=8'hE3;
    mem['h1C20]=8'h73; mem['h1C21]=8'h23; mem['h1C22]=8'h72; mem['h1C23]=8'hE1;
    mem['h1C24]=8'hC9; mem['h1C25]=8'hCD; mem['h1C26]=8'h50; mem['h1C27]=8'h0D;
    mem['h1C28]=8'hCD; mem['h1C29]=8'h92; mem['h1C2A]=8'h09; mem['h1C2B]=8'hC5;
    mem['h1C2C]=8'h21; mem['h1C2D]=8'h2E; mem['h1C2E]=8'h81; mem['h1C2F]=8'h7A;
    mem['h1C30]=8'hFE; mem['h1C31]=8'h00; mem['h1C32]=8'h28; mem['h1C33]=8'h0C;
    mem['h1C34]=8'hCD; mem['h1C35]=8'h5D; mem['h1C36]=8'h1C; mem['h1C37]=8'h78;
    mem['h1C38]=8'hFE; mem['h1C39]=8'h30; mem['h1C3A]=8'h28; mem['h1C3B]=8'h02;
    mem['h1C3C]=8'h70; mem['h1C3D]=8'h23; mem['h1C3E]=8'h71; mem['h1C3F]=8'h23;
    mem['h1C40]=8'h7B; mem['h1C41]=8'hCD; mem['h1C42]=8'h5D; mem['h1C43]=8'h1C;
    mem['h1C44]=8'h7A; mem['h1C45]=8'hFE; mem['h1C46]=8'h00; mem['h1C47]=8'h20;
    mem['h1C48]=8'h05; mem['h1C49]=8'h78; mem['h1C4A]=8'hFE; mem['h1C4B]=8'h30;
    mem['h1C4C]=8'h28; mem['h1C4D]=8'h02; mem['h1C4E]=8'h70; mem['h1C4F]=8'h23;
    mem['h1C50]=8'h71; mem['h1C51]=8'h23; mem['h1C52]=8'hAF; mem['h1C53]=8'h77;
    mem['h1C54]=8'h23; mem['h1C55]=8'h77; mem['h1C56]=8'hC1; mem['h1C57]=8'h21;
    mem['h1C58]=8'h2E; mem['h1C59]=8'h81; mem['h1C5A]=8'hC3; mem['h1C5B]=8'hB6;
    mem['h1C5C]=8'h11; mem['h1C5D]=8'h47; mem['h1C5E]=8'hE6; mem['h1C5F]=8'h0F;
    mem['h1C60]=8'hFE; mem['h1C61]=8'h0A; mem['h1C62]=8'h38; mem['h1C63]=8'h02;
    mem['h1C64]=8'hC6; mem['h1C65]=8'h07; mem['h1C66]=8'hC6; mem['h1C67]=8'h30;
    mem['h1C68]=8'h4F; mem['h1C69]=8'h78; mem['h1C6A]=8'h0F; mem['h1C6B]=8'h0F;
    mem['h1C6C]=8'h0F; mem['h1C6D]=8'h0F; mem['h1C6E]=8'hE6; mem['h1C6F]=8'h0F;
    mem['h1C70]=8'hFE; mem['h1C71]=8'h0A; mem['h1C72]=8'h38; mem['h1C73]=8'h02;
    mem['h1C74]=8'hC6; mem['h1C75]=8'h07; mem['h1C76]=8'hC6; mem['h1C77]=8'h30;
    mem['h1C78]=8'h47; mem['h1C79]=8'hC9; mem['h1C7A]=8'hEB; mem['h1C7B]=8'h21;
    mem['h1C7C]=8'h00; mem['h1C7D]=8'h00; mem['h1C7E]=8'hCD; mem['h1C7F]=8'h93;
    mem['h1C80]=8'h1C; mem['h1C81]=8'hDA; mem['h1C82]=8'hB3; mem['h1C83]=8'h1C;
    mem['h1C84]=8'h18; mem['h1C85]=8'h05; mem['h1C86]=8'hCD; mem['h1C87]=8'h93;
    mem['h1C88]=8'h1C; mem['h1C89]=8'h38; mem['h1C8A]=8'h1F; mem['h1C8B]=8'h29;
    mem['h1C8C]=8'h29; mem['h1C8D]=8'h29; mem['h1C8E]=8'h29; mem['h1C8F]=8'hB5;
    mem['h1C90]=8'h6F; mem['h1C91]=8'h18; mem['h1C92]=8'hF3; mem['h1C93]=8'h13;
    mem['h1C94]=8'h1A; mem['h1C95]=8'hFE; mem['h1C96]=8'h20; mem['h1C97]=8'hCA;
    mem['h1C98]=8'h93; mem['h1C99]=8'h1C; mem['h1C9A]=8'hD6; mem['h1C9B]=8'h30;
    mem['h1C9C]=8'hD8; mem['h1C9D]=8'hFE; mem['h1C9E]=8'h0A; mem['h1C9F]=8'h38;
    mem['h1CA0]=8'h05; mem['h1CA1]=8'hD6; mem['h1CA2]=8'h07; mem['h1CA3]=8'hFE;
    mem['h1CA4]=8'h0A; mem['h1CA5]=8'hD8; mem['h1CA6]=8'hFE; mem['h1CA7]=8'h10;
    mem['h1CA8]=8'h3F; mem['h1CA9]=8'hC9; mem['h1CAA]=8'hEB; mem['h1CAB]=8'h7A;
    mem['h1CAC]=8'h4B; mem['h1CAD]=8'hE5; mem['h1CAE]=8'hCD; mem['h1CAF]=8'h07;
    mem['h1CB0]=8'h11; mem['h1CB1]=8'hE1; mem['h1CB2]=8'hC9; mem['h1CB3]=8'h1E;
    mem['h1CB4]=8'h26; mem['h1CB5]=8'hC3; mem['h1CB6]=8'h9C; mem['h1CB7]=8'h04;
    mem['h1CB8]=8'hCD; mem['h1CB9]=8'h50; mem['h1CBA]=8'h0D; mem['h1CBB]=8'hCD;
    mem['h1CBC]=8'h92; mem['h1CBD]=8'h09; mem['h1CBE]=8'hC5; mem['h1CBF]=8'h21;
    mem['h1CC0]=8'h2E; mem['h1CC1]=8'h81; mem['h1CC2]=8'h06; mem['h1CC3]=8'h11;
    mem['h1CC4]=8'h05; mem['h1CC5]=8'h78; mem['h1CC6]=8'hFE; mem['h1CC7]=8'h01;
    mem['h1CC8]=8'h28; mem['h1CC9]=8'h08; mem['h1CCA]=8'hCB; mem['h1CCB]=8'h13;
    mem['h1CCC]=8'hCB; mem['h1CCD]=8'h12; mem['h1CCE]=8'h30; mem['h1CCF]=8'hF4;
    mem['h1CD0]=8'h18; mem['h1CD1]=8'h04; mem['h1CD2]=8'hCB; mem['h1CD3]=8'h13;
    mem['h1CD4]=8'hCB; mem['h1CD5]=8'h12; mem['h1CD6]=8'h3E; mem['h1CD7]=8'h30;
    mem['h1CD8]=8'hCE; mem['h1CD9]=8'h00; mem['h1CDA]=8'h77; mem['h1CDB]=8'h23;
    mem['h1CDC]=8'h05; mem['h1CDD]=8'h20; mem['h1CDE]=8'hF3; mem['h1CDF]=8'hAF;
    mem['h1CE0]=8'h77; mem['h1CE1]=8'h23; mem['h1CE2]=8'h77; mem['h1CE3]=8'hC1;
    mem['h1CE4]=8'h21; mem['h1CE5]=8'h2E; mem['h1CE6]=8'h81; mem['h1CE7]=8'hC3;
    mem['h1CE8]=8'hB6; mem['h1CE9]=8'h11; mem['h1CEA]=8'hEB; mem['h1CEB]=8'h21;
    mem['h1CEC]=8'h00; mem['h1CED]=8'h00; mem['h1CEE]=8'hCD; mem['h1CEF]=8'h07;
    mem['h1CF0]=8'h1D; mem['h1CF1]=8'hDA; mem['h1CF2]=8'h15; mem['h1CF3]=8'h1D;
    mem['h1CF4]=8'hD6; mem['h1CF5]=8'h30; mem['h1CF6]=8'h29; mem['h1CF7]=8'hB5;
    mem['h1CF8]=8'h6F; mem['h1CF9]=8'hCD; mem['h1CFA]=8'h07; mem['h1CFB]=8'h1D;
    mem['h1CFC]=8'h30; mem['h1CFD]=8'hF6; mem['h1CFE]=8'hEB; mem['h1CFF]=8'h7A;
    mem['h1D00]=8'h4B; mem['h1D01]=8'hE5; mem['h1D02]=8'hCD; mem['h1D03]=8'h07;
    mem['h1D04]=8'h11; mem['h1D05]=8'hE1; mem['h1D06]=8'hC9; mem['h1D07]=8'h13;
    mem['h1D08]=8'h1A; mem['h1D09]=8'hFE; mem['h1D0A]=8'h20; mem['h1D0B]=8'hCA;
    mem['h1D0C]=8'h07; mem['h1D0D]=8'h1D; mem['h1D0E]=8'hFE; mem['h1D0F]=8'h30;
    mem['h1D10]=8'hD8; mem['h1D11]=8'hFE; mem['h1D12]=8'h32; mem['h1D13]=8'h3F;
    mem['h1D14]=8'hC9; mem['h1D15]=8'h1E; mem['h1D16]=8'h28; mem['h1D17]=8'hC3;
    mem['h1D18]=8'h9C; mem['h1D19]=8'h04; mem['h1D1A]=8'hC3; mem['h1D1B]=8'hE1;
    mem['h1D1C]=8'h00; mem['h1D1D]=8'hC3; mem['h1D1E]=8'h08; mem['h1D1F]=8'h00;
    mem['h1D20]=8'hC3; mem['h1D21]=8'h00; mem['h1D22]=8'h00; mem['h1D23]=8'h3E;
    mem['h1D24]=8'h00; mem['h1D25]=8'h32; mem['h1D26]=8'h92; mem['h1D27]=8'h80;
    mem['h1D28]=8'hC3; mem['h1D29]=8'hE8; mem['h1D2A]=8'h00; mem['h1D2B]=8'hF5;
    mem['h1D2C]=8'hA0; mem['h1D2D]=8'hC1; mem['h1D2E]=8'hB8; mem['h1D2F]=8'h3E;
    mem['h1D30]=8'h00; mem['h1D31]=8'hC9; mem['h1D32]=8'hCD; mem['h1D33]=8'h61;
    mem['h1D34]=8'h07; mem['h1D35]=8'hC3; mem['h1D36]=8'h88; mem['h1D37]=8'h0B;
    mem['h1D38]=8'hFF; mem['h1D39]=8'hFF; mem['h1D3A]=8'hFF; mem['h1D3B]=8'hFF;
    mem['h1D3C]=8'hFF; mem['h1D3D]=8'hFF; mem['h1D3E]=8'hFF; mem['h1D3F]=8'hFF;
    mem['h1D40]=8'hFF; mem['h1D41]=8'hFF; mem['h1D42]=8'hFF; mem['h1D43]=8'hFF;
    mem['h1D44]=8'hFF; mem['h1D45]=8'hFF; mem['h1D46]=8'hFF; mem['h1D47]=8'hFF;
    mem['h1D48]=8'hFF; mem['h1D49]=8'hFF; mem['h1D4A]=8'hFF; mem['h1D4B]=8'hFF;
    mem['h1D4C]=8'hFF; mem['h1D4D]=8'hFF; mem['h1D4E]=8'hFF; mem['h1D4F]=8'hFF;
    mem['h1D50]=8'hFF; mem['h1D51]=8'hFF; mem['h1D52]=8'hFF; mem['h1D53]=8'hFF;
    mem['h1D54]=8'hFF; mem['h1D55]=8'hFF; mem['h1D56]=8'hFF; mem['h1D57]=8'hFF;
    mem['h1D58]=8'hFF; mem['h1D59]=8'hFF; mem['h1D5A]=8'hFF; mem['h1D5B]=8'hFF;
    mem['h1D5C]=8'hFF; mem['h1D5D]=8'hFF; mem['h1D5E]=8'hFF; mem['h1D5F]=8'hFF;
    mem['h1D60]=8'hFF; mem['h1D61]=8'hFF; mem['h1D62]=8'hFF; mem['h1D63]=8'hFF;
    mem['h1D64]=8'hFF; mem['h1D65]=8'hFF; mem['h1D66]=8'hFF; mem['h1D67]=8'hFF;
    mem['h1D68]=8'hFF; mem['h1D69]=8'hFF; mem['h1D6A]=8'hFF; mem['h1D6B]=8'hFF;
    mem['h1D6C]=8'hFF; mem['h1D6D]=8'hFF; mem['h1D6E]=8'hFF; mem['h1D6F]=8'hFF;
    mem['h1D70]=8'hFF; mem['h1D71]=8'hFF; mem['h1D72]=8'hFF; mem['h1D73]=8'hFF;
    mem['h1D74]=8'hFF; mem['h1D75]=8'hFF; mem['h1D76]=8'hFF; mem['h1D77]=8'hFF;
    mem['h1D78]=8'hFF; mem['h1D79]=8'hFF; mem['h1D7A]=8'hFF; mem['h1D7B]=8'hFF;
    mem['h1D7C]=8'hFF; mem['h1D7D]=8'hFF; mem['h1D7E]=8'hFF; mem['h1D7F]=8'hFF;
    mem['h1D80]=8'hFF; mem['h1D81]=8'hFF; mem['h1D82]=8'hFF; mem['h1D83]=8'hFF;
    mem['h1D84]=8'hFF; mem['h1D85]=8'hFF; mem['h1D86]=8'hFF; mem['h1D87]=8'hFF;
    mem['h1D88]=8'hFF; mem['h1D89]=8'hFF; mem['h1D8A]=8'hFF; mem['h1D8B]=8'hFF;
    mem['h1D8C]=8'hFF; mem['h1D8D]=8'hFF; mem['h1D8E]=8'hFF; mem['h1D8F]=8'hFF;
    mem['h1D90]=8'hFF; mem['h1D91]=8'hFF; mem['h1D92]=8'hFF; mem['h1D93]=8'hFF;
    mem['h1D94]=8'hFF; mem['h1D95]=8'hFF; mem['h1D96]=8'hFF; mem['h1D97]=8'hFF;
    mem['h1D98]=8'hFF; mem['h1D99]=8'hFF; mem['h1D9A]=8'hFF; mem['h1D9B]=8'hFF;
    mem['h1D9C]=8'hFF; mem['h1D9D]=8'hFF; mem['h1D9E]=8'hFF; mem['h1D9F]=8'hFF;
    mem['h1DA0]=8'hFF; mem['h1DA1]=8'hFF; mem['h1DA2]=8'hFF; mem['h1DA3]=8'hFF;
    mem['h1DA4]=8'hFF; mem['h1DA5]=8'hFF; mem['h1DA6]=8'hFF; mem['h1DA7]=8'hFF;
    mem['h1DA8]=8'hFF; mem['h1DA9]=8'hFF; mem['h1DAA]=8'hFF; mem['h1DAB]=8'hFF;
    mem['h1DAC]=8'hFF; mem['h1DAD]=8'hFF; mem['h1DAE]=8'hFF; mem['h1DAF]=8'hFF;
    mem['h1DB0]=8'hFF; mem['h1DB1]=8'hFF; mem['h1DB2]=8'hFF; mem['h1DB3]=8'hFF;
    mem['h1DB4]=8'hFF; mem['h1DB5]=8'hFF; mem['h1DB6]=8'hFF; mem['h1DB7]=8'hFF;
    mem['h1DB8]=8'hFF; mem['h1DB9]=8'hFF; mem['h1DBA]=8'hFF; mem['h1DBB]=8'hFF;
    mem['h1DBC]=8'hFF; mem['h1DBD]=8'hFF; mem['h1DBE]=8'hFF; mem['h1DBF]=8'hFF;
    mem['h1DC0]=8'hFF; mem['h1DC1]=8'hFF; mem['h1DC2]=8'hFF; mem['h1DC3]=8'hFF;
    mem['h1DC4]=8'hFF; mem['h1DC5]=8'hFF; mem['h1DC6]=8'hFF; mem['h1DC7]=8'hFF;
    mem['h1DC8]=8'hFF; mem['h1DC9]=8'hFF; mem['h1DCA]=8'hFF; mem['h1DCB]=8'hFF;
    mem['h1DCC]=8'hFF; mem['h1DCD]=8'hFF; mem['h1DCE]=8'hFF; mem['h1DCF]=8'hFF;
    mem['h1DD0]=8'hFF; mem['h1DD1]=8'hFF; mem['h1DD2]=8'hFF; mem['h1DD3]=8'hFF;
    mem['h1DD4]=8'hFF; mem['h1DD5]=8'hFF; mem['h1DD6]=8'hFF; mem['h1DD7]=8'hFF;
    mem['h1DD8]=8'hFF; mem['h1DD9]=8'hFF; mem['h1DDA]=8'hFF; mem['h1DDB]=8'hFF;
    mem['h1DDC]=8'hFF; mem['h1DDD]=8'hFF; mem['h1DDE]=8'hFF; mem['h1DDF]=8'hFF;
    mem['h1DE0]=8'hFF; mem['h1DE1]=8'hFF; mem['h1DE2]=8'hFF; mem['h1DE3]=8'hFF;
    mem['h1DE4]=8'hFF; mem['h1DE5]=8'hFF; mem['h1DE6]=8'hFF; mem['h1DE7]=8'hFF;
    mem['h1DE8]=8'hFF; mem['h1DE9]=8'hFF; mem['h1DEA]=8'hFF; mem['h1DEB]=8'hFF;
    mem['h1DEC]=8'hFF; mem['h1DED]=8'hFF; mem['h1DEE]=8'hFF; mem['h1DEF]=8'hFF;
    mem['h1DF0]=8'hFF; mem['h1DF1]=8'hFF; mem['h1DF2]=8'hFF; mem['h1DF3]=8'hFF;
    mem['h1DF4]=8'hFF; mem['h1DF5]=8'hFF; mem['h1DF6]=8'hFF; mem['h1DF7]=8'hFF;
    mem['h1DF8]=8'hFF; mem['h1DF9]=8'hFF; mem['h1DFA]=8'hFF; mem['h1DFB]=8'hFF;
    mem['h1DFC]=8'hFF; mem['h1DFD]=8'hFF; mem['h1DFE]=8'hFF; mem['h1DFF]=8'hFF;
    mem['h1E00]=8'hFF; mem['h1E01]=8'hFF; mem['h1E02]=8'hFF; mem['h1E03]=8'hFF;
    mem['h1E04]=8'hFF; mem['h1E05]=8'hFF; mem['h1E06]=8'hFF; mem['h1E07]=8'hFF;
    mem['h1E08]=8'hFF; mem['h1E09]=8'hFF; mem['h1E0A]=8'hFF; mem['h1E0B]=8'hFF;
    mem['h1E0C]=8'hFF; mem['h1E0D]=8'hFF; mem['h1E0E]=8'hFF; mem['h1E0F]=8'hFF;
    mem['h1E10]=8'hFF; mem['h1E11]=8'hFF; mem['h1E12]=8'hFF; mem['h1E13]=8'hFF;
    mem['h1E14]=8'hFF; mem['h1E15]=8'hFF; mem['h1E16]=8'hFF; mem['h1E17]=8'hFF;
    mem['h1E18]=8'hFF; mem['h1E19]=8'hFF; mem['h1E1A]=8'hFF; mem['h1E1B]=8'hFF;
    mem['h1E1C]=8'hFF; mem['h1E1D]=8'hFF; mem['h1E1E]=8'hFF; mem['h1E1F]=8'hFF;
    mem['h1E20]=8'hFF; mem['h1E21]=8'hFF; mem['h1E22]=8'hFF; mem['h1E23]=8'hFF;
    mem['h1E24]=8'hFF; mem['h1E25]=8'hFF; mem['h1E26]=8'hFF; mem['h1E27]=8'hFF;
    mem['h1E28]=8'hFF; mem['h1E29]=8'hFF; mem['h1E2A]=8'hFF; mem['h1E2B]=8'hFF;
    mem['h1E2C]=8'hFF; mem['h1E2D]=8'hFF; mem['h1E2E]=8'hFF; mem['h1E2F]=8'hFF;
    mem['h1E30]=8'hFF; mem['h1E31]=8'hFF; mem['h1E32]=8'hFF; mem['h1E33]=8'hFF;
    mem['h1E34]=8'hFF; mem['h1E35]=8'hFF; mem['h1E36]=8'hFF; mem['h1E37]=8'hFF;
    mem['h1E38]=8'hFF; mem['h1E39]=8'hFF; mem['h1E3A]=8'hFF; mem['h1E3B]=8'hFF;
    mem['h1E3C]=8'hFF; mem['h1E3D]=8'hFF; mem['h1E3E]=8'hFF; mem['h1E3F]=8'hFF;
    mem['h1E40]=8'hFF; mem['h1E41]=8'hFF; mem['h1E42]=8'hFF; mem['h1E43]=8'hFF;
    mem['h1E44]=8'hFF; mem['h1E45]=8'hFF; mem['h1E46]=8'hFF; mem['h1E47]=8'hFF;
    mem['h1E48]=8'hFF; mem['h1E49]=8'hFF; mem['h1E4A]=8'hFF; mem['h1E4B]=8'hFF;
    mem['h1E4C]=8'hFF; mem['h1E4D]=8'hFF; mem['h1E4E]=8'hFF; mem['h1E4F]=8'hFF;
    mem['h1E50]=8'hFF; mem['h1E51]=8'hFF; mem['h1E52]=8'hFF; mem['h1E53]=8'hFF;
    mem['h1E54]=8'hFF; mem['h1E55]=8'hFF; mem['h1E56]=8'hFF; mem['h1E57]=8'hFF;
    mem['h1E58]=8'hFF; mem['h1E59]=8'hFF; mem['h1E5A]=8'hFF; mem['h1E5B]=8'hFF;
    mem['h1E5C]=8'hFF; mem['h1E5D]=8'hFF; mem['h1E5E]=8'hFF; mem['h1E5F]=8'hFF;
    mem['h1E60]=8'hFF; mem['h1E61]=8'hFF; mem['h1E62]=8'hFF; mem['h1E63]=8'hFF;
    mem['h1E64]=8'hFF; mem['h1E65]=8'hFF; mem['h1E66]=8'hFF; mem['h1E67]=8'hFF;
    mem['h1E68]=8'hFF; mem['h1E69]=8'hFF; mem['h1E6A]=8'hFF; mem['h1E6B]=8'hFF;
    mem['h1E6C]=8'hFF; mem['h1E6D]=8'hFF; mem['h1E6E]=8'hFF; mem['h1E6F]=8'hFF;
    mem['h1E70]=8'hFF; mem['h1E71]=8'hFF; mem['h1E72]=8'hFF; mem['h1E73]=8'hFF;
    mem['h1E74]=8'hFF; mem['h1E75]=8'hFF; mem['h1E76]=8'hFF; mem['h1E77]=8'hFF;
    mem['h1E78]=8'hFF; mem['h1E79]=8'hFF; mem['h1E7A]=8'hFF; mem['h1E7B]=8'hFF;
    mem['h1E7C]=8'hFF; mem['h1E7D]=8'hFF; mem['h1E7E]=8'hFF; mem['h1E7F]=8'hFF;
    mem['h1E80]=8'hFF; mem['h1E81]=8'hFF; mem['h1E82]=8'hFF; mem['h1E83]=8'hFF;
    mem['h1E84]=8'hFF; mem['h1E85]=8'hFF; mem['h1E86]=8'hFF; mem['h1E87]=8'hFF;
    mem['h1E88]=8'hFF; mem['h1E89]=8'hFF; mem['h1E8A]=8'hFF; mem['h1E8B]=8'hFF;
    mem['h1E8C]=8'hFF; mem['h1E8D]=8'hFF; mem['h1E8E]=8'hFF; mem['h1E8F]=8'hFF;
    mem['h1E90]=8'hFF; mem['h1E91]=8'hFF; mem['h1E92]=8'hFF; mem['h1E93]=8'hFF;
    mem['h1E94]=8'hFF; mem['h1E95]=8'hFF; mem['h1E96]=8'hFF; mem['h1E97]=8'hFF;
    mem['h1E98]=8'hFF; mem['h1E99]=8'hFF; mem['h1E9A]=8'hFF; mem['h1E9B]=8'hFF;
    mem['h1E9C]=8'hFF; mem['h1E9D]=8'hFF; mem['h1E9E]=8'hFF; mem['h1E9F]=8'hFF;
    mem['h1EA0]=8'hFF; mem['h1EA1]=8'hFF; mem['h1EA2]=8'hFF; mem['h1EA3]=8'hFF;
    mem['h1EA4]=8'hFF; mem['h1EA5]=8'hFF; mem['h1EA6]=8'hFF; mem['h1EA7]=8'hFF;
    mem['h1EA8]=8'hFF; mem['h1EA9]=8'hFF; mem['h1EAA]=8'hFF; mem['h1EAB]=8'hFF;
    mem['h1EAC]=8'hFF; mem['h1EAD]=8'hFF; mem['h1EAE]=8'hFF; mem['h1EAF]=8'hFF;
    mem['h1EB0]=8'hFF; mem['h1EB1]=8'hFF; mem['h1EB2]=8'hFF; mem['h1EB3]=8'hFF;
    mem['h1EB4]=8'hFF; mem['h1EB5]=8'hFF; mem['h1EB6]=8'hFF; mem['h1EB7]=8'hFF;
    mem['h1EB8]=8'hFF; mem['h1EB9]=8'hFF; mem['h1EBA]=8'hFF; mem['h1EBB]=8'hFF;
    mem['h1EBC]=8'hFF; mem['h1EBD]=8'hFF; mem['h1EBE]=8'hFF; mem['h1EBF]=8'hFF;
    mem['h1EC0]=8'hFF; mem['h1EC1]=8'hFF; mem['h1EC2]=8'hFF; mem['h1EC3]=8'hFF;
    mem['h1EC4]=8'hFF; mem['h1EC5]=8'hFF; mem['h1EC6]=8'hFF; mem['h1EC7]=8'hFF;
    mem['h1EC8]=8'hFF; mem['h1EC9]=8'hFF; mem['h1ECA]=8'hFF; mem['h1ECB]=8'hFF;
    mem['h1ECC]=8'hFF; mem['h1ECD]=8'hFF; mem['h1ECE]=8'hFF; mem['h1ECF]=8'hFF;
    mem['h1ED0]=8'hFF; mem['h1ED1]=8'hFF; mem['h1ED2]=8'hFF; mem['h1ED3]=8'hFF;
    mem['h1ED4]=8'hFF; mem['h1ED5]=8'hFF; mem['h1ED6]=8'hFF; mem['h1ED7]=8'hFF;
    mem['h1ED8]=8'hFF; mem['h1ED9]=8'hFF; mem['h1EDA]=8'hFF; mem['h1EDB]=8'hFF;
    mem['h1EDC]=8'hFF; mem['h1EDD]=8'hFF; mem['h1EDE]=8'hFF; mem['h1EDF]=8'hFF;
    mem['h1EE0]=8'hFF; mem['h1EE1]=8'hFF; mem['h1EE2]=8'hFF; mem['h1EE3]=8'hFF;
    mem['h1EE4]=8'hFF; mem['h1EE5]=8'hFF; mem['h1EE6]=8'hFF; mem['h1EE7]=8'hFF;
    mem['h1EE8]=8'hFF; mem['h1EE9]=8'hFF; mem['h1EEA]=8'hFF; mem['h1EEB]=8'hFF;
    mem['h1EEC]=8'hFF; mem['h1EED]=8'hFF; mem['h1EEE]=8'hFF; mem['h1EEF]=8'hFF;
    mem['h1EF0]=8'hFF; mem['h1EF1]=8'hFF; mem['h1EF2]=8'hFF; mem['h1EF3]=8'hFF;
    mem['h1EF4]=8'hFF; mem['h1EF5]=8'hFF; mem['h1EF6]=8'hFF; mem['h1EF7]=8'hFF;
    mem['h1EF8]=8'hFF; mem['h1EF9]=8'hFF; mem['h1EFA]=8'hFF; mem['h1EFB]=8'hFF;
    mem['h1EFC]=8'hFF; mem['h1EFD]=8'hFF; mem['h1EFE]=8'hFF; mem['h1EFF]=8'hFF;
    mem['h1F00]=8'hFF; mem['h1F01]=8'hFF; mem['h1F02]=8'hFF; mem['h1F03]=8'hFF;
    mem['h1F04]=8'hFF; mem['h1F05]=8'hFF; mem['h1F06]=8'hFF; mem['h1F07]=8'hFF;
    mem['h1F08]=8'hFF; mem['h1F09]=8'hFF; mem['h1F0A]=8'hFF; mem['h1F0B]=8'hFF;
    mem['h1F0C]=8'hFF; mem['h1F0D]=8'hFF; mem['h1F0E]=8'hFF; mem['h1F0F]=8'hFF;
    mem['h1F10]=8'hFF; mem['h1F11]=8'hFF; mem['h1F12]=8'hFF; mem['h1F13]=8'hFF;
    mem['h1F14]=8'hFF; mem['h1F15]=8'hFF; mem['h1F16]=8'hFF; mem['h1F17]=8'hFF;
    mem['h1F18]=8'hFF; mem['h1F19]=8'hFF; mem['h1F1A]=8'hFF; mem['h1F1B]=8'hFF;
    mem['h1F1C]=8'hFF; mem['h1F1D]=8'hFF; mem['h1F1E]=8'hFF; mem['h1F1F]=8'hFF;
    mem['h1F20]=8'hFF; mem['h1F21]=8'hFF; mem['h1F22]=8'hFF; mem['h1F23]=8'hFF;
    mem['h1F24]=8'hFF; mem['h1F25]=8'hFF; mem['h1F26]=8'hFF; mem['h1F27]=8'hFF;
    mem['h1F28]=8'hFF; mem['h1F29]=8'hFF; mem['h1F2A]=8'hFF; mem['h1F2B]=8'hFF;
    mem['h1F2C]=8'hFF; mem['h1F2D]=8'hFF; mem['h1F2E]=8'hFF; mem['h1F2F]=8'hFF;
    mem['h1F30]=8'hFF; mem['h1F31]=8'hFF; mem['h1F32]=8'hFF; mem['h1F33]=8'hFF;
    mem['h1F34]=8'hFF; mem['h1F35]=8'hFF; mem['h1F36]=8'hFF; mem['h1F37]=8'hFF;
    mem['h1F38]=8'hFF; mem['h1F39]=8'hFF; mem['h1F3A]=8'hFF; mem['h1F3B]=8'hFF;
    mem['h1F3C]=8'hFF; mem['h1F3D]=8'hFF; mem['h1F3E]=8'hFF; mem['h1F3F]=8'hFF;
    mem['h1F40]=8'hFF; mem['h1F41]=8'hFF; mem['h1F42]=8'hFF; mem['h1F43]=8'hFF;
    mem['h1F44]=8'hFF; mem['h1F45]=8'hFF; mem['h1F46]=8'hFF; mem['h1F47]=8'hFF;
    mem['h1F48]=8'hFF; mem['h1F49]=8'hFF; mem['h1F4A]=8'hFF; mem['h1F4B]=8'hFF;
    mem['h1F4C]=8'hFF; mem['h1F4D]=8'hFF; mem['h1F4E]=8'hFF; mem['h1F4F]=8'hFF;
    mem['h1F50]=8'hFF; mem['h1F51]=8'hFF; mem['h1F52]=8'hFF; mem['h1F53]=8'hFF;
    mem['h1F54]=8'hFF; mem['h1F55]=8'hFF; mem['h1F56]=8'hFF; mem['h1F57]=8'hFF;
    mem['h1F58]=8'hFF; mem['h1F59]=8'hFF; mem['h1F5A]=8'hFF; mem['h1F5B]=8'hFF;
    mem['h1F5C]=8'hFF; mem['h1F5D]=8'hFF; mem['h1F5E]=8'hFF; mem['h1F5F]=8'hFF;
    mem['h1F60]=8'hFF; mem['h1F61]=8'hFF; mem['h1F62]=8'hFF; mem['h1F63]=8'hFF;
    mem['h1F64]=8'hFF; mem['h1F65]=8'hFF; mem['h1F66]=8'hFF; mem['h1F67]=8'hFF;
    mem['h1F68]=8'hFF; mem['h1F69]=8'hFF; mem['h1F6A]=8'hFF; mem['h1F6B]=8'hFF;
    mem['h1F6C]=8'hFF; mem['h1F6D]=8'hFF; mem['h1F6E]=8'hFF; mem['h1F6F]=8'hFF;
    mem['h1F70]=8'hFF; mem['h1F71]=8'hFF; mem['h1F72]=8'hFF; mem['h1F73]=8'hFF;
    mem['h1F74]=8'hFF; mem['h1F75]=8'hFF; mem['h1F76]=8'hFF; mem['h1F77]=8'hFF;
    mem['h1F78]=8'hFF; mem['h1F79]=8'hFF; mem['h1F7A]=8'hFF; mem['h1F7B]=8'hFF;
    mem['h1F7C]=8'hFF; mem['h1F7D]=8'hFF; mem['h1F7E]=8'hFF; mem['h1F7F]=8'hFF;
    mem['h1F80]=8'hFF; mem['h1F81]=8'hFF; mem['h1F82]=8'hFF; mem['h1F83]=8'hFF;
    mem['h1F84]=8'hFF; mem['h1F85]=8'hFF; mem['h1F86]=8'hFF; mem['h1F87]=8'hFF;
    mem['h1F88]=8'hFF; mem['h1F89]=8'hFF; mem['h1F8A]=8'hFF; mem['h1F8B]=8'hFF;
    mem['h1F8C]=8'hFF; mem['h1F8D]=8'hFF; mem['h1F8E]=8'hFF; mem['h1F8F]=8'hFF;
    mem['h1F90]=8'hFF; mem['h1F91]=8'hFF; mem['h1F92]=8'hFF; mem['h1F93]=8'hFF;
    mem['h1F94]=8'hFF; mem['h1F95]=8'hFF; mem['h1F96]=8'hFF; mem['h1F97]=8'hFF;
    mem['h1F98]=8'hFF; mem['h1F99]=8'hFF; mem['h1F9A]=8'hFF; mem['h1F9B]=8'hFF;
    mem['h1F9C]=8'hFF; mem['h1F9D]=8'hFF; mem['h1F9E]=8'hFF; mem['h1F9F]=8'hFF;
    mem['h1FA0]=8'hFF; mem['h1FA1]=8'hFF; mem['h1FA2]=8'hFF; mem['h1FA3]=8'hFF;
    mem['h1FA4]=8'hFF; mem['h1FA5]=8'hFF; mem['h1FA6]=8'hFF; mem['h1FA7]=8'hFF;
    mem['h1FA8]=8'hFF; mem['h1FA9]=8'hFF; mem['h1FAA]=8'hFF; mem['h1FAB]=8'hFF;
    mem['h1FAC]=8'hFF; mem['h1FAD]=8'hFF; mem['h1FAE]=8'hFF; mem['h1FAF]=8'hFF;
    mem['h1FB0]=8'hFF; mem['h1FB1]=8'hFF; mem['h1FB2]=8'hFF; mem['h1FB3]=8'hFF;
    mem['h1FB4]=8'hFF; mem['h1FB5]=8'hFF; mem['h1FB6]=8'hFF; mem['h1FB7]=8'hFF;
    mem['h1FB8]=8'hFF; mem['h1FB9]=8'hFF; mem['h1FBA]=8'hFF; mem['h1FBB]=8'hFF;
    mem['h1FBC]=8'hFF; mem['h1FBD]=8'hFF; mem['h1FBE]=8'hFF; mem['h1FBF]=8'hFF;
    mem['h1FC0]=8'hFF; mem['h1FC1]=8'hFF; mem['h1FC2]=8'hFF; mem['h1FC3]=8'hFF;
    mem['h1FC4]=8'hFF; mem['h1FC5]=8'hFF; mem['h1FC6]=8'hFF; mem['h1FC7]=8'hFF;
    mem['h1FC8]=8'hFF; mem['h1FC9]=8'hFF; mem['h1FCA]=8'hFF; mem['h1FCB]=8'hFF;
    mem['h1FCC]=8'hFF; mem['h1FCD]=8'hFF; mem['h1FCE]=8'hFF; mem['h1FCF]=8'hFF;
    mem['h1FD0]=8'hFF; mem['h1FD1]=8'hFF; mem['h1FD2]=8'hFF; mem['h1FD3]=8'hFF;
    mem['h1FD4]=8'hFF; mem['h1FD5]=8'hFF; mem['h1FD6]=8'hFF; mem['h1FD7]=8'hFF;
    mem['h1FD8]=8'hFF; mem['h1FD9]=8'hFF; mem['h1FDA]=8'hFF; mem['h1FDB]=8'hFF;
    mem['h1FDC]=8'hFF; mem['h1FDD]=8'hFF; mem['h1FDE]=8'hFF; mem['h1FDF]=8'hFF;
    mem['h1FE0]=8'hFF; mem['h1FE1]=8'hFF; mem['h1FE2]=8'hFF; mem['h1FE3]=8'hFF;
    mem['h1FE4]=8'hFF; mem['h1FE5]=8'hFF; mem['h1FE6]=8'hFF; mem['h1FE7]=8'hFF;
    mem['h1FE8]=8'hFF; mem['h1FE9]=8'hFF; mem['h1FEA]=8'hFF; mem['h1FEB]=8'hFF;
    mem['h1FEC]=8'hFF; mem['h1FED]=8'hFF; mem['h1FEE]=8'hFF; mem['h1FEF]=8'hFF;
    mem['h1FF0]=8'hFF; mem['h1FF1]=8'hFF; mem['h1FF2]=8'hFF; mem['h1FF3]=8'hFF;
    mem['h1FF4]=8'hFF; mem['h1FF5]=8'hFF; mem['h1FF6]=8'hFF; mem['h1FF7]=8'hFF;
    mem['h1FF8]=8'hFF; mem['h1FF9]=8'hFF; mem['h1FFA]=8'hFF; mem['h1FFB]=8'hFF;
    mem['h1FFC]=8'hFF; mem['h1FFD]=8'hFF; mem['h1FFE]=8'hFF; mem['h1FFF]=8'hFF;
end
