// rom.v
// to be included from the top module at the compile

initial
begin
    mem['h0000]=8'hC0; mem['h0001]=8'h44; mem['h0002]=8'h00; mem['h0003]=8'h01;
    mem['h0004]=8'hFF; mem['h0005]=8'hFF; mem['h0006]=8'hFF; mem['h0007]=8'hFF;
    mem['h0008]=8'h44; mem['h0009]=8'h00; mem['h000A]=8'h01; mem['h000B]=8'hFF;
    mem['h000C]=8'hFF; mem['h000D]=8'hFF; mem['h000E]=8'hFF; mem['h000F]=8'hFF;
    mem['h0010]=8'h44; mem['h0011]=8'h00; mem['h0012]=8'h01; mem['h0013]=8'hFF;
    mem['h0014]=8'hFF; mem['h0015]=8'hFF; mem['h0016]=8'hFF; mem['h0017]=8'hFF;
    mem['h0018]=8'h44; mem['h0019]=8'h00; mem['h001A]=8'h01; mem['h001B]=8'hFF;
    mem['h001C]=8'hFF; mem['h001D]=8'hFF; mem['h001E]=8'hFF; mem['h001F]=8'hFF;
    mem['h0020]=8'h44; mem['h0021]=8'h00; mem['h0022]=8'h01; mem['h0023]=8'hFF;
    mem['h0024]=8'hFF; mem['h0025]=8'hFF; mem['h0026]=8'hFF; mem['h0027]=8'hFF;
    mem['h0028]=8'h44; mem['h0029]=8'h00; mem['h002A]=8'h01; mem['h002B]=8'hFF;
    mem['h002C]=8'hFF; mem['h002D]=8'hFF; mem['h002E]=8'hFF; mem['h002F]=8'hFF;
    mem['h0030]=8'h44; mem['h0031]=8'h00; mem['h0032]=8'h01; mem['h0033]=8'hFF;
    mem['h0034]=8'hFF; mem['h0035]=8'hFF; mem['h0036]=8'hFF; mem['h0037]=8'hFF;
    mem['h0038]=8'h44; mem['h0039]=8'h00; mem['h003A]=8'h01; mem['h003B]=8'hFF;
    mem['h003C]=8'hFF; mem['h003D]=8'hFF; mem['h003E]=8'hFF; mem['h003F]=8'hFF;
    mem['h0040]=8'hC8; mem['h0041]=8'h41; mem['h0042]=8'h24; mem['h0043]=8'h04;
    mem['h0044]=8'h68; mem['h0045]=8'h41; mem['h0046]=8'h00; mem['h0047]=8'hC1;
    mem['h0048]=8'h61; mem['h0049]=8'h07; mem['h004A]=8'h41; mem['h004B]=8'h24;
    mem['h004C]=8'h01; mem['h004D]=8'h68; mem['h004E]=8'h4A; mem['h004F]=8'h00;
    mem['h0050]=8'h43; mem['h0051]=8'h07; mem['h0052]=8'hC7; mem['h0053]=8'hA0;
    mem['h0054]=8'h2B; mem['h0055]=8'h46; mem['h0056]=8'h40; mem['h0057]=8'h00;
    mem['h0058]=8'h30; mem['h0059]=8'h48; mem['h005A]=8'h52; mem['h005B]=8'h00;
    mem['h005C]=8'h28; mem['h005D]=8'h44; mem['h005E]=8'h52; mem['h005F]=8'h00;
    mem['h0060]=8'h06; mem['h0061]=8'h0D; mem['h0062]=8'h46; mem['h0063]=8'h40;
    mem['h0064]=8'h00; mem['h0065]=8'h06; mem['h0066]=8'h0A; mem['h0067]=8'h46;
    mem['h0068]=8'h40; mem['h0069]=8'h00; mem['h006A]=8'h07; mem['h006B]=8'hFF;
    mem['h006C]=8'hFF; mem['h006D]=8'hFF; mem['h006E]=8'hFF; mem['h006F]=8'hFF;
    mem['h0070]=8'hFF; mem['h0071]=8'hFF; mem['h0072]=8'hFF; mem['h0073]=8'hFF;
    mem['h0074]=8'hFF; mem['h0075]=8'hFF; mem['h0076]=8'hFF; mem['h0077]=8'hFF;
    mem['h0078]=8'hFF; mem['h0079]=8'hFF; mem['h007A]=8'hFF; mem['h007B]=8'hFF;
    mem['h007C]=8'hFF; mem['h007D]=8'hFF; mem['h007E]=8'hFF; mem['h007F]=8'hFF;
    mem['h0080]=8'hFF; mem['h0081]=8'hFF; mem['h0082]=8'hFF; mem['h0083]=8'hFF;
    mem['h0084]=8'hFF; mem['h0085]=8'hFF; mem['h0086]=8'hFF; mem['h0087]=8'hFF;
    mem['h0088]=8'hFF; mem['h0089]=8'hFF; mem['h008A]=8'hFF; mem['h008B]=8'hFF;
    mem['h008C]=8'hFF; mem['h008D]=8'hFF; mem['h008E]=8'hFF; mem['h008F]=8'hFF;
    mem['h0090]=8'hFF; mem['h0091]=8'hFF; mem['h0092]=8'hFF; mem['h0093]=8'hFF;
    mem['h0094]=8'hFF; mem['h0095]=8'hFF; mem['h0096]=8'hFF; mem['h0097]=8'hFF;
    mem['h0098]=8'hFF; mem['h0099]=8'hFF; mem['h009A]=8'hFF; mem['h009B]=8'hFF;
    mem['h009C]=8'hFF; mem['h009D]=8'hFF; mem['h009E]=8'hFF; mem['h009F]=8'hFF;
    mem['h00A0]=8'hFF; mem['h00A1]=8'hFF; mem['h00A2]=8'hFF; mem['h00A3]=8'hFF;
    mem['h00A4]=8'hFF; mem['h00A5]=8'hFF; mem['h00A6]=8'hFF; mem['h00A7]=8'hFF;
    mem['h00A8]=8'hFF; mem['h00A9]=8'hFF; mem['h00AA]=8'hFF; mem['h00AB]=8'hFF;
    mem['h00AC]=8'hFF; mem['h00AD]=8'hFF; mem['h00AE]=8'hFF; mem['h00AF]=8'hFF;
    mem['h00B0]=8'hFF; mem['h00B1]=8'hFF; mem['h00B2]=8'hFF; mem['h00B3]=8'hFF;
    mem['h00B4]=8'hFF; mem['h00B5]=8'hFF; mem['h00B6]=8'hFF; mem['h00B7]=8'hFF;
    mem['h00B8]=8'hFF; mem['h00B9]=8'hFF; mem['h00BA]=8'hFF; mem['h00BB]=8'hFF;
    mem['h00BC]=8'hFF; mem['h00BD]=8'hFF; mem['h00BE]=8'hFF; mem['h00BF]=8'hFF;
    mem['h00C0]=8'hFF; mem['h00C1]=8'hFF; mem['h00C2]=8'hFF; mem['h00C3]=8'hFF;
    mem['h00C4]=8'hFF; mem['h00C5]=8'hFF; mem['h00C6]=8'hFF; mem['h00C7]=8'hFF;
    mem['h00C8]=8'hFF; mem['h00C9]=8'hFF; mem['h00CA]=8'hFF; mem['h00CB]=8'hFF;
    mem['h00CC]=8'hFF; mem['h00CD]=8'hFF; mem['h00CE]=8'hFF; mem['h00CF]=8'hFF;
    mem['h00D0]=8'hFF; mem['h00D1]=8'hFF; mem['h00D2]=8'hFF; mem['h00D3]=8'hFF;
    mem['h00D4]=8'hFF; mem['h00D5]=8'hFF; mem['h00D6]=8'hFF; mem['h00D7]=8'hFF;
    mem['h00D8]=8'hFF; mem['h00D9]=8'hFF; mem['h00DA]=8'hFF; mem['h00DB]=8'hFF;
    mem['h00DC]=8'hFF; mem['h00DD]=8'hFF; mem['h00DE]=8'hFF; mem['h00DF]=8'hFF;
    mem['h00E0]=8'hFF; mem['h00E1]=8'hFF; mem['h00E2]=8'hFF; mem['h00E3]=8'hFF;
    mem['h00E4]=8'hFF; mem['h00E5]=8'hFF; mem['h00E6]=8'hFF; mem['h00E7]=8'hFF;
    mem['h00E8]=8'hFF; mem['h00E9]=8'hFF; mem['h00EA]=8'hFF; mem['h00EB]=8'hFF;
    mem['h00EC]=8'hFF; mem['h00ED]=8'hFF; mem['h00EE]=8'hFF; mem['h00EF]=8'hFF;
    mem['h00F0]=8'hFF; mem['h00F1]=8'hFF; mem['h00F2]=8'hFF; mem['h00F3]=8'hFF;
    mem['h00F4]=8'hFF; mem['h00F5]=8'hFF; mem['h00F6]=8'hFF; mem['h00F7]=8'hFF;
    mem['h00F8]=8'hFF; mem['h00F9]=8'hFF; mem['h00FA]=8'hFF; mem['h00FB]=8'hFF;
    mem['h00FC]=8'hFF; mem['h00FD]=8'hFF; mem['h00FE]=8'hFF; mem['h00FF]=8'hFF;
    mem['h0100]=8'h2E; mem['h0101]=8'h01; mem['h0102]=8'h36; mem['h0103]=8'h0A;
    mem['h0104]=8'h46; mem['h0105]=8'h52; mem['h0106]=8'h00; mem['h0107]=8'h44;
    mem['h0108]=8'h89; mem['h0109]=8'h07; mem['h010A]=8'h1B; mem['h010B]=8'h40;
    mem['h010C]=8'h1F; mem['h010D]=8'h02; mem['h010E]=8'h00; mem['h010F]=8'h0D;
    mem['h0110]=8'h0A; mem['h0111]=8'h56; mem['h0112]=8'h54; mem['h0113]=8'h4C;
    mem['h0114]=8'h2D; mem['h0115]=8'h38; mem['h0116]=8'h30; mem['h0117]=8'h30;
    mem['h0118]=8'h38; mem['h0119]=8'h20; mem['h011A]=8'h49; mem['h011B]=8'h6E;
    mem['h011C]=8'h74; mem['h011D]=8'h65; mem['h011E]=8'h72; mem['h011F]=8'h70;
    mem['h0120]=8'h72; mem['h0121]=8'h65; mem['h0122]=8'h74; mem['h0123]=8'h65;
    mem['h0124]=8'h72; mem['h0125]=8'h20; mem['h0126]=8'h56; mem['h0127]=8'h65;
    mem['h0128]=8'h72; mem['h0129]=8'h20; mem['h012A]=8'h32; mem['h012B]=8'h2E;
    mem['h012C]=8'h30; mem['h012D]=8'h0D; mem['h012E]=8'h0A; mem['h012F]=8'h28;
    mem['h0130]=8'h43; mem['h0131]=8'h29; mem['h0132]=8'h20; mem['h0133]=8'h32;
    mem['h0134]=8'h30; mem['h0135]=8'h32; mem['h0136]=8'h34; mem['h0137]=8'h20;
    mem['h0138]=8'h52; mem['h0139]=8'h79; mem['h013A]=8'h6F; mem['h013B]=8'h20;
    mem['h013C]=8'h4D; mem['h013D]=8'h75; mem['h013E]=8'h6B; mem['h013F]=8'h61;
    mem['h0140]=8'h69; mem['h0141]=8'h0D; mem['h0142]=8'h0A; mem['h0143]=8'h00;
    mem['h0144]=8'h0D; mem['h0145]=8'h0A; mem['h0146]=8'h4F; mem['h0147]=8'h4B;
    mem['h0148]=8'h0D; mem['h0149]=8'h0A; mem['h014A]=8'h00; mem['h014B]=8'h53;
    mem['h014C]=8'h59; mem['h014D]=8'h45; mem['h014E]=8'h52; mem['h014F]=8'h52;
    mem['h0150]=8'h00; mem['h0151]=8'h50; mem['h0152]=8'h52; mem['h0153]=8'h45;
    mem['h0154]=8'h52; mem['h0155]=8'h52; mem['h0156]=8'h00; mem['h0157]=8'h4F;
    mem['h0158]=8'h50; mem['h0159]=8'h45; mem['h015A]=8'h52; mem['h015B]=8'h52;
    mem['h015C]=8'h00; mem['h015D]=8'h45; mem['h015E]=8'h4F; mem['h015F]=8'h4C;
    mem['h0160]=8'h45; mem['h0161]=8'h52; mem['h0162]=8'h52; mem['h0163]=8'h00;
    mem['h0164]=8'h46; mem['h0165]=8'h54; mem['h0166]=8'h45; mem['h0167]=8'h52;
    mem['h0168]=8'h52; mem['h0169]=8'h00; mem['h016A]=8'h42; mem['h016B]=8'h55;
    mem['h016C]=8'h46; mem['h016D]=8'h3D; mem['h016E]=8'h00; mem['h016F]=8'h53;
    mem['h0170]=8'h50; mem['h0171]=8'h3D; mem['h0172]=8'h00; mem['h0173]=8'h50;
    mem['h0174]=8'h43; mem['h0175]=8'h53; mem['h0176]=8'h50; mem['h0177]=8'h3D;
    mem['h0178]=8'h00; mem['h0179]=8'h49; mem['h017A]=8'h4E; mem['h017B]=8'h20;
    mem['h017C]=8'h23; mem['h017D]=8'h00; mem['h017E]=8'h2E; mem['h017F]=8'h3E;
    mem['h0180]=8'h36; mem['h0181]=8'h00; mem['h0182]=8'hF7; mem['h0183]=8'h31;
    mem['h0184]=8'hF9; mem['h0185]=8'h31; mem['h0186]=8'hFA; mem['h0187]=8'hD6;
    mem['h0188]=8'h36; mem['h0189]=8'h00; mem['h018A]=8'hFA; mem['h018B]=8'hF2;
    mem['h018C]=8'hD7; mem['h018D]=8'h07; mem['h018E]=8'h46; mem['h018F]=8'hCE;
    mem['h0190]=8'h01; mem['h0191]=8'h2E; mem['h0192]=8'h3E; mem['h0193]=8'h36;
    mem['h0194]=8'h00; mem['h0195]=8'hF7; mem['h0196]=8'hD7; mem['h0197]=8'h30;
    mem['h0198]=8'h30; mem['h0199]=8'hCE; mem['h019A]=8'h36; mem['h019B]=8'h00;
    mem['h019C]=8'hF9; mem['h019D]=8'hF1; mem['h019E]=8'h31; mem['h019F]=8'hCF;
    mem['h01A0]=8'h2E; mem['h01A1]=8'h38; mem['h01A2]=8'h36; mem['h01A3]=8'h7C;
    mem['h01A4]=8'h3E; mem['h01A5]=8'h44; mem['h01A6]=8'h30; mem['h01A7]=8'hFA;
    mem['h01A8]=8'h30; mem['h01A9]=8'hF9; mem['h01AA]=8'h46; mem['h01AB]=8'h0C;
    mem['h01AC]=8'h02; mem['h01AD]=8'h44; mem['h01AE]=8'h7C; mem['h01AF]=8'h38;
    mem['h01B0]=8'h2E; mem['h01B1]=8'h3F; mem['h01B2]=8'h36; mem['h01B3]=8'h00;
    mem['h01B4]=8'hF7; mem['h01B5]=8'h31; mem['h01B6]=8'hF8; mem['h01B7]=8'hC6;
    mem['h01B8]=8'h36; mem['h01B9]=8'h00; mem['h01BA]=8'hF8; mem['h01BB]=8'hF7;
    mem['h01BC]=8'hC7; mem['h01BD]=8'h07; mem['h01BE]=8'h2E; mem['h01BF]=8'h3F;
    mem['h01C0]=8'h36; mem['h01C1]=8'h00; mem['h01C2]=8'hF7; mem['h01C3]=8'h31;
    mem['h01C4]=8'hF8; mem['h01C5]=8'h31; mem['h01C6]=8'hF9; mem['h01C7]=8'hCE;
    mem['h01C8]=8'h36; mem['h01C9]=8'h00; mem['h01CA]=8'hF9; mem['h01CB]=8'hF1;
    mem['h01CC]=8'hCF; mem['h01CD]=8'h07; mem['h01CE]=8'h2E; mem['h01CF]=8'h3F;
    mem['h01D0]=8'h36; mem['h01D1]=8'h00; mem['h01D2]=8'hF7; mem['h01D3]=8'h31;
    mem['h01D4]=8'hF9; mem['h01D5]=8'h31; mem['h01D6]=8'hFA; mem['h01D7]=8'hD6;
    mem['h01D8]=8'h36; mem['h01D9]=8'h00; mem['h01DA]=8'hFA; mem['h01DB]=8'hF2;
    mem['h01DC]=8'hD7; mem['h01DD]=8'h07; mem['h01DE]=8'h2E; mem['h01DF]=8'h3F;
    mem['h01E0]=8'h36; mem['h01E1]=8'h00; mem['h01E2]=8'hF7; mem['h01E3]=8'h31;
    mem['h01E4]=8'hFB; mem['h01E5]=8'h31; mem['h01E6]=8'hFC; mem['h01E7]=8'hE6;
    mem['h01E8]=8'h36; mem['h01E9]=8'h00; mem['h01EA]=8'hFC; mem['h01EB]=8'hF4;
    mem['h01EC]=8'hE7; mem['h01ED]=8'h07; mem['h01EE]=8'h2E; mem['h01EF]=8'h3F;
    mem['h01F0]=8'h36; mem['h01F1]=8'h00; mem['h01F2]=8'hF7; mem['h01F3]=8'h30;
    mem['h01F4]=8'hC6; mem['h01F5]=8'h36; mem['h01F6]=8'h00; mem['h01F7]=8'hF8;
    mem['h01F8]=8'hF0; mem['h01F9]=8'h31; mem['h01FA]=8'hC7; mem['h01FB]=8'h07;
    mem['h01FC]=8'h2E; mem['h01FD]=8'h3F; mem['h01FE]=8'h36; mem['h01FF]=8'h00;
    mem['h0200]=8'hF7; mem['h0201]=8'hCF; mem['h0202]=8'h30; mem['h0203]=8'h30;
    mem['h0204]=8'hC6; mem['h0205]=8'h36; mem['h0206]=8'h00; mem['h0207]=8'hF8;
    mem['h0208]=8'hF0; mem['h0209]=8'h31; mem['h020A]=8'hC7; mem['h020B]=8'h07;
    mem['h020C]=8'h2E; mem['h020D]=8'h3F; mem['h020E]=8'h36; mem['h020F]=8'h00;
    mem['h0210]=8'hF7; mem['h0211]=8'hD7; mem['h0212]=8'h30; mem['h0213]=8'h30;
    mem['h0214]=8'hCE; mem['h0215]=8'h36; mem['h0216]=8'h00; mem['h0217]=8'hF9;
    mem['h0218]=8'hF1; mem['h0219]=8'h31; mem['h021A]=8'hCF; mem['h021B]=8'h07;
    mem['h021C]=8'h2E; mem['h021D]=8'h3F; mem['h021E]=8'h36; mem['h021F]=8'h00;
    mem['h0220]=8'hF7; mem['h0221]=8'hE7; mem['h0222]=8'h30; mem['h0223]=8'h30;
    mem['h0224]=8'hDE; mem['h0225]=8'h36; mem['h0226]=8'h00; mem['h0227]=8'hFB;
    mem['h0228]=8'hF3; mem['h0229]=8'h31; mem['h022A]=8'hDF; mem['h022B]=8'h07;
    mem['h022C]=8'h2E; mem['h022D]=8'h38; mem['h022E]=8'h36; mem['h022F]=8'h5C;
    mem['h0230]=8'hFA; mem['h0231]=8'h30; mem['h0232]=8'hF9; mem['h0233]=8'hF0;
    mem['h0234]=8'hD7; mem['h0235]=8'h30; mem['h0236]=8'hCF; mem['h0237]=8'h46;
    mem['h0238]=8'hCE; mem['h0239]=8'h01; mem['h023A]=8'h2E; mem['h023B]=8'h38;
    mem['h023C]=8'h36; mem['h023D]=8'h5C; mem['h023E]=8'hD7; mem['h023F]=8'h30;
    mem['h0240]=8'hCF; mem['h0241]=8'h07; mem['h0242]=8'h2E; mem['h0243]=8'h38;
    mem['h0244]=8'h36; mem['h0245]=8'h5C; mem['h0246]=8'hFA; mem['h0247]=8'h30;
    mem['h0248]=8'hF9; mem['h0249]=8'h46; mem['h024A]=8'h0C; mem['h024B]=8'h02;
    mem['h024C]=8'h2E; mem['h024D]=8'h38; mem['h024E]=8'hF0; mem['h024F]=8'hFA;
    mem['h0250]=8'h30; mem['h0251]=8'hF9; mem['h0252]=8'h36; mem['h0253]=8'h5C;
    mem['h0254]=8'hD7; mem['h0255]=8'h30; mem['h0256]=8'hCF; mem['h0257]=8'h07;
    mem['h0258]=8'h2E; mem['h0259]=8'h38; mem['h025A]=8'hF4; mem['h025B]=8'hC7;
    mem['h025C]=8'hF3; mem['h025D]=8'hF8; mem['h025E]=8'hF4; mem['h025F]=8'h30;
    mem['h0260]=8'hC7; mem['h0261]=8'hF3; mem['h0262]=8'h30; mem['h0263]=8'hF8;
    mem['h0264]=8'h07; mem['h0265]=8'h2E; mem['h0266]=8'h38; mem['h0267]=8'hF3;
    mem['h0268]=8'hC7; mem['h0269]=8'hF4; mem['h026A]=8'hF8; mem['h026B]=8'hF3;
    mem['h026C]=8'h30; mem['h026D]=8'hC7; mem['h026E]=8'hF4; mem['h026F]=8'h30;
    mem['h0270]=8'hF8; mem['h0271]=8'h07; mem['h0272]=8'h2E; mem['h0273]=8'h38;
    mem['h0274]=8'hF3; mem['h0275]=8'hC7; mem['h0276]=8'hF1; mem['h0277]=8'hF8;
    mem['h0278]=8'hF3; mem['h0279]=8'h30; mem['h027A]=8'hC7; mem['h027B]=8'hF1;
    mem['h027C]=8'h30; mem['h027D]=8'hF8; mem['h027E]=8'h07; mem['h027F]=8'h2E;
    mem['h0280]=8'h38; mem['h0281]=8'hF1; mem['h0282]=8'hC7; mem['h0283]=8'hF3;
    mem['h0284]=8'hF8; mem['h0285]=8'hF1; mem['h0286]=8'h30; mem['h0287]=8'hC7;
    mem['h0288]=8'hF3; mem['h0289]=8'h30; mem['h028A]=8'hF8; mem['h028B]=8'h07;
    mem['h028C]=8'h2E; mem['h028D]=8'h38; mem['h028E]=8'hF4; mem['h028F]=8'hC7;
    mem['h0290]=8'hF1; mem['h0291]=8'hF8; mem['h0292]=8'hF4; mem['h0293]=8'h30;
    mem['h0294]=8'hC7; mem['h0295]=8'hF1; mem['h0296]=8'h30; mem['h0297]=8'hF8;
    mem['h0298]=8'h07; mem['h0299]=8'h2E; mem['h029A]=8'h38; mem['h029B]=8'hF3;
    mem['h029C]=8'hCF; mem['h029D]=8'h08; mem['h029E]=8'hF9; mem['h029F]=8'h0B;
    mem['h02A0]=8'h30; mem['h02A1]=8'hCF; mem['h02A2]=8'h08; mem['h02A3]=8'hF9;
    mem['h02A4]=8'h07; mem['h02A5]=8'h2E; mem['h02A6]=8'h38; mem['h02A7]=8'hF3;
    mem['h02A8]=8'hCF; mem['h02A9]=8'h08; mem['h02AA]=8'h09; mem['h02AB]=8'h68;
    mem['h02AC]=8'hB1; mem['h02AD]=8'h02; mem['h02AE]=8'h09; mem['h02AF]=8'hF9;
    mem['h02B0]=8'h07; mem['h02B1]=8'h09; mem['h02B2]=8'hF9; mem['h02B3]=8'h30;
    mem['h02B4]=8'hCF; mem['h02B5]=8'h09; mem['h02B6]=8'hF9; mem['h02B7]=8'h07;
    mem['h02B8]=8'h46; mem['h02B9]=8'hBE; mem['h02BA]=8'h01; mem['h02BB]=8'hF0;
    mem['h02BC]=8'h0A; mem['h02BD]=8'h0A; mem['h02BE]=8'h0A; mem['h02BF]=8'h0A;
    mem['h02C0]=8'h24; mem['h02C1]=8'h0F; mem['h02C2]=8'h3C; mem['h02C3]=8'h0A;
    mem['h02C4]=8'h60; mem['h02C5]=8'hC9; mem['h02C6]=8'h02; mem['h02C7]=8'h04;
    mem['h02C8]=8'h07; mem['h02C9]=8'h04; mem['h02CA]=8'h30; mem['h02CB]=8'h46;
    mem['h02CC]=8'h40; mem['h02CD]=8'h00; mem['h02CE]=8'hC6; mem['h02CF]=8'h24;
    mem['h02D0]=8'h0F; mem['h02D1]=8'h3C; mem['h02D2]=8'h0A; mem['h02D3]=8'h60;
    mem['h02D4]=8'hD8; mem['h02D5]=8'h02; mem['h02D6]=8'h04; mem['h02D7]=8'h07;
    mem['h02D8]=8'h04; mem['h02D9]=8'h30; mem['h02DA]=8'h46; mem['h02DB]=8'h40;
    mem['h02DC]=8'h00; mem['h02DD]=8'h44; mem['h02DE]=8'hFC; mem['h02DF]=8'h01;
    mem['h02E0]=8'h3C; mem['h02E1]=8'h30; mem['h02E2]=8'h60; mem['h02E3]=8'hE8;
    mem['h02E4]=8'h02; mem['h02E5]=8'h3C; mem['h02E6]=8'h3A; mem['h02E7]=8'h07;
    mem['h02E8]=8'hA0; mem['h02E9]=8'h07; mem['h02EA]=8'h3C; mem['h02EB]=8'h30;
    mem['h02EC]=8'h60; mem['h02ED]=8'h02; mem['h02EE]=8'h03; mem['h02EF]=8'h3C;
    mem['h02F0]=8'h3A; mem['h02F1]=8'h23; mem['h02F2]=8'h3C; mem['h02F3]=8'h41;
    mem['h02F4]=8'h60; mem['h02F5]=8'h02; mem['h02F6]=8'h03; mem['h02F7]=8'h3C;
    mem['h02F8]=8'h47; mem['h02F9]=8'h23; mem['h02FA]=8'h3C; mem['h02FB]=8'h61;
    mem['h02FC]=8'h60; mem['h02FD]=8'h02; mem['h02FE]=8'h03; mem['h02FF]=8'h3C;
    mem['h0300]=8'h67; mem['h0301]=8'h23; mem['h0302]=8'hA0; mem['h0303]=8'h07;
    mem['h0304]=8'h3C; mem['h0305]=8'h41; mem['h0306]=8'h60; mem['h0307]=8'h14;
    mem['h0308]=8'h03; mem['h0309]=8'h3C; mem['h030A]=8'h5B; mem['h030B]=8'h23;
    mem['h030C]=8'h3C; mem['h030D]=8'h61; mem['h030E]=8'h60; mem['h030F]=8'h14;
    mem['h0310]=8'h03; mem['h0311]=8'h3C; mem['h0312]=8'h7B; mem['h0313]=8'h23;
    mem['h0314]=8'hA0; mem['h0315]=8'h07; mem['h0316]=8'h14; mem['h0317]=8'h30;
    mem['h0318]=8'h3C; mem['h0319]=8'h0A; mem['h031A]=8'h23; mem['h031B]=8'h24;
    mem['h031C]=8'h1F; mem['h031D]=8'h14; mem['h031E]=8'h07; mem['h031F]=8'h07;
    mem['h0320]=8'h46; mem['h0321]=8'hCE; mem['h0322]=8'h01; mem['h0323]=8'h2E;
    mem['h0324]=8'h38; mem['h0325]=8'hF3; mem['h0326]=8'hD7; mem['h0327]=8'h30;
    mem['h0328]=8'hCF; mem['h0329]=8'hE9; mem['h032A]=8'hF2; mem['h032B]=8'hC7;
    mem['h032C]=8'h44; mem['h032D]=8'h0C; mem['h032E]=8'h02; mem['h032F]=8'h46;
    mem['h0330]=8'hCE; mem['h0331]=8'h01; mem['h0332]=8'h2E; mem['h0333]=8'h38;
    mem['h0334]=8'hF3; mem['h0335]=8'hD7; mem['h0336]=8'h30; mem['h0337]=8'hCF;
    mem['h0338]=8'hE9; mem['h0339]=8'hF2; mem['h033A]=8'hF8; mem['h033B]=8'h44;
    mem['h033C]=8'h0C; mem['h033D]=8'h02; mem['h033E]=8'h46; mem['h033F]=8'hDE;
    mem['h0340]=8'h01; mem['h0341]=8'h2E; mem['h0342]=8'h38; mem['h0343]=8'hF3;
    mem['h0344]=8'hE7; mem['h0345]=8'h30; mem['h0346]=8'hDF; mem['h0347]=8'hEB;
    mem['h0348]=8'hF4; mem['h0349]=8'hD7; mem['h034A]=8'h30; mem['h034B]=8'h48;
    mem['h034C]=8'h4F; mem['h034D]=8'h03; mem['h034E]=8'h28; mem['h034F]=8'hCF;
    mem['h0350]=8'h44; mem['h0351]=8'h1C; mem['h0352]=8'h02; mem['h0353]=8'h46;
    mem['h0354]=8'hDE; mem['h0355]=8'h01; mem['h0356]=8'h2E; mem['h0357]=8'h38;
    mem['h0358]=8'hF3; mem['h0359]=8'hE7; mem['h035A]=8'h30; mem['h035B]=8'hDF;
    mem['h035C]=8'hEB; mem['h035D]=8'hF4; mem['h035E]=8'hFA; mem['h035F]=8'h30;
    mem['h0360]=8'h48; mem['h0361]=8'h64; mem['h0362]=8'h03; mem['h0363]=8'h28;
    mem['h0364]=8'hF9; mem['h0365]=8'h44; mem['h0366]=8'h1C; mem['h0367]=8'h02;
    mem['h0368]=8'h46; mem['h0369]=8'hCE; mem['h036A]=8'h01; mem['h036B]=8'h46;
    mem['h036C]=8'hDE; mem['h036D]=8'h01; mem['h036E]=8'h2E; mem['h036F]=8'h38;
    mem['h0370]=8'hF3; mem['h0371]=8'hE7; mem['h0372]=8'h30; mem['h0373]=8'hDF;
    mem['h0374]=8'hEB; mem['h0375]=8'hF4; mem['h0376]=8'hD7; mem['h0377]=8'h30;
    mem['h0378]=8'h48; mem['h0379]=8'h7C; mem['h037A]=8'h03; mem['h037B]=8'h28;
    mem['h037C]=8'hCF; mem['h037D]=8'h46; mem['h037E]=8'h1C; mem['h037F]=8'h02;
    mem['h0380]=8'h2E; mem['h0381]=8'h38; mem['h0382]=8'hF4; mem['h0383]=8'hFA;
    mem['h0384]=8'h30; mem['h0385]=8'hF9; mem['h0386]=8'h44; mem['h0387]=8'h0C;
    mem['h0388]=8'h02; mem['h0389]=8'h46; mem['h038A]=8'hCE; mem['h038B]=8'h01;
    mem['h038C]=8'h46; mem['h038D]=8'hDE; mem['h038E]=8'h01; mem['h038F]=8'h2E;
    mem['h0390]=8'h38; mem['h0391]=8'hF4; mem['h0392]=8'hD7; mem['h0393]=8'h30;
    mem['h0394]=8'hCF; mem['h0395]=8'hF3; mem['h0396]=8'hE7; mem['h0397]=8'h30;
    mem['h0398]=8'hDF; mem['h0399]=8'hEB; mem['h039A]=8'hF4; mem['h039B]=8'hFA;
    mem['h039C]=8'h30; mem['h039D]=8'h48; mem['h039E]=8'hA1; mem['h039F]=8'h03;
    mem['h03A0]=8'h28; mem['h03A1]=8'hF9; mem['h03A2]=8'h46; mem['h03A3]=8'h1C;
    mem['h03A4]=8'h02; mem['h03A5]=8'h44; mem['h03A6]=8'h0C; mem['h03A7]=8'h02;
    mem['h03A8]=8'h46; mem['h03A9]=8'hCE; mem['h03AA]=8'h01; mem['h03AB]=8'h46;
    mem['h03AC]=8'hDE; mem['h03AD]=8'h01; mem['h03AE]=8'h26; mem['h03AF]=8'h52;
    mem['h03B0]=8'h46; mem['h03B1]=8'h65; mem['h03B2]=8'h02; mem['h03B3]=8'h46;
    mem['h03B4]=8'h4A; mem['h03B5]=8'h00; mem['h03B6]=8'h3C; mem['h03B7]=8'h0D;
    mem['h03B8]=8'h48; mem['h03B9]=8'hC1; mem['h03BA]=8'h03; mem['h03BB]=8'h46;
    mem['h03BC]=8'h60; mem['h03BD]=8'h00; mem['h03BE]=8'h44; mem['h03BF]=8'hF2;
    mem['h03C0]=8'h03; mem['h03C1]=8'h3C; mem['h03C2]=8'h08; mem['h03C3]=8'h48;
    mem['h03C4]=8'hE6; mem['h03C5]=8'h03; mem['h03C6]=8'h26; mem['h03C7]=8'h52;
    mem['h03C8]=8'h46; mem['h03C9]=8'hFC; mem['h03CA]=8'h06; mem['h03CB]=8'h48;
    mem['h03CC]=8'hD1; mem['h03CD]=8'h03; mem['h03CE]=8'h44; mem['h03CF]=8'hB3;
    mem['h03D0]=8'h03; mem['h03D1]=8'h46; mem['h03D2]=8'hA5; mem['h03D3]=8'h02;
    mem['h03D4]=8'h06; mem['h03D5]=8'h08; mem['h03D6]=8'h46; mem['h03D7]=8'h40;
    mem['h03D8]=8'h00; mem['h03D9]=8'h06; mem['h03DA]=8'h20; mem['h03DB]=8'h46;
    mem['h03DC]=8'h40; mem['h03DD]=8'h00; mem['h03DE]=8'h06; mem['h03DF]=8'h08;
    mem['h03E0]=8'h46; mem['h03E1]=8'h40; mem['h03E2]=8'h00; mem['h03E3]=8'h44;
    mem['h03E4]=8'hB3; mem['h03E5]=8'h03; mem['h03E6]=8'h46; mem['h03E7]=8'h40;
    mem['h03E8]=8'h00; mem['h03E9]=8'h46; mem['h03EA]=8'h2F; mem['h03EB]=8'h03;
    mem['h03EC]=8'h46; mem['h03ED]=8'h99; mem['h03EE]=8'h02; mem['h03EF]=8'h44;
    mem['h03F0]=8'hB3; mem['h03F1]=8'h03; mem['h03F2]=8'hA8; mem['h03F3]=8'h46;
    mem['h03F4]=8'h2F; mem['h03F5]=8'h03; mem['h03F6]=8'h46; mem['h03F7]=8'h99;
    mem['h03F8]=8'h02; mem['h03F9]=8'h46; mem['h03FA]=8'h2F; mem['h03FB]=8'h03;
    mem['h03FC]=8'h46; mem['h03FD]=8'h58; mem['h03FE]=8'h02; mem['h03FF]=8'h46;
    mem['h0400]=8'h1C; mem['h0401]=8'h02; mem['h0402]=8'h44; mem['h0403]=8'h0C;
    mem['h0404]=8'h02; mem['h0405]=8'h46; mem['h0406]=8'hBE; mem['h0407]=8'h01;
    mem['h0408]=8'h46; mem['h0409]=8'h12; mem['h040A]=8'h05; mem['h040B]=8'h46;
    mem['h040C]=8'h20; mem['h040D]=8'h03; mem['h040E]=8'h46; mem['h040F]=8'hEA;
    mem['h0410]=8'h02; mem['h0411]=8'h40; mem['h0412]=8'h2E; mem['h0413]=8'h04;
    mem['h0414]=8'h46; mem['h0415]=8'h99; mem['h0416]=8'h02; mem['h0417]=8'h46;
    mem['h0418]=8'h16; mem['h0419]=8'h03; mem['h041A]=8'hC8; mem['h041B]=8'hC4;
    mem['h041C]=8'h46; mem['h041D]=8'h99; mem['h041E]=8'h05; mem['h041F]=8'h46;
    mem['h0420]=8'h99; mem['h0421]=8'h05; mem['h0422]=8'h46; mem['h0423]=8'h99;
    mem['h0424]=8'h05; mem['h0425]=8'h46; mem['h0426]=8'h99; mem['h0427]=8'h05;
    mem['h0428]=8'h46; mem['h0429]=8'h61; mem['h042A]=8'h05; mem['h042B]=8'h44;
    mem['h042C]=8'h0B; mem['h042D]=8'h04; mem['h042E]=8'h44; mem['h042F]=8'hFC;
    mem['h0430]=8'h01; mem['h0431]=8'h46; mem['h0432]=8'h20; mem['h0433]=8'h03;
    mem['h0434]=8'h3C; mem['h0435]=8'h30; mem['h0436]=8'h68; mem['h0437]=8'h05;
    mem['h0438]=8'h04; mem['h0439]=8'h46; mem['h043A]=8'hB0; mem['h043B]=8'h01;
    mem['h043C]=8'h46; mem['h043D]=8'hCE; mem['h043E]=8'h01; mem['h043F]=8'h46;
    mem['h0440]=8'h12; mem['h0441]=8'h05; mem['h0442]=8'hD3; mem['h0443]=8'hDA;
    mem['h0444]=8'hC2; mem['h0445]=8'h46; mem['h0446]=8'h20; mem['h0447]=8'h03;
    mem['h0448]=8'h46; mem['h0449]=8'hE0; mem['h044A]=8'h02; mem['h044B]=8'h40;
    mem['h044C]=8'h74; mem['h044D]=8'h04; mem['h044E]=8'h46; mem['h044F]=8'h99;
    mem['h0450]=8'h02; mem['h0451]=8'h46; mem['h0452]=8'h16; mem['h0453]=8'h03;
    mem['h0454]=8'hC8; mem['h0455]=8'hC4; mem['h0456]=8'h46; mem['h0457]=8'h99;
    mem['h0458]=8'h05; mem['h0459]=8'h1E; mem['h045A]=8'h5A; mem['h045B]=8'h46;
    mem['h045C]=8'h58; mem['h045D]=8'h02; mem['h045E]=8'hC4; mem['h045F]=8'h46;
    mem['h0460]=8'h99; mem['h0461]=8'h05; mem['h0462]=8'h46; mem['h0463]=8'h99;
    mem['h0464]=8'h05; mem['h0465]=8'h1E; mem['h0466]=8'h5A; mem['h0467]=8'h46;
    mem['h0468]=8'h6D; mem['h0469]=8'h05; mem['h046A]=8'hC3; mem['h046B]=8'h46;
    mem['h046C]=8'h61; mem['h046D]=8'h05; mem['h046E]=8'h46; mem['h046F]=8'h65;
    mem['h0470]=8'h02; mem['h0471]=8'h44; mem['h0472]=8'h43; mem['h0473]=8'h04;
    mem['h0474]=8'h46; mem['h0475]=8'h0C; mem['h0476]=8'h02; mem['h0477]=8'h44;
    mem['h0478]=8'hEE; mem['h0479]=8'h01; mem['h047A]=8'h46; mem['h047B]=8'h99;
    mem['h047C]=8'h02; mem['h047D]=8'h46; mem['h047E]=8'h20; mem['h047F]=8'h03;
    mem['h0480]=8'h3C; mem['h0481]=8'h63; mem['h0482]=8'h68; mem['h0483]=8'h8D;
    mem['h0484]=8'h04; mem['h0485]=8'h3C; mem['h0486]=8'h64; mem['h0487]=8'h68;
    mem['h0488]=8'hAF; mem['h0489]=8'h04; mem['h048A]=8'h44; mem['h048B]=8'hD8;
    mem['h048C]=8'h07; mem['h048D]=8'h46; mem['h048E]=8'hCE; mem['h048F]=8'h01;
    mem['h0490]=8'h2E; mem['h0491]=8'h10; mem['h0492]=8'h36; mem['h0493]=8'h00;
    mem['h0494]=8'h0E; mem['h0495]=8'h37; mem['h0496]=8'h16; mem['h0497]=8'hFF;
    mem['h0498]=8'h3E; mem['h0499]=8'h00; mem['h049A]=8'h30; mem['h049B]=8'h48;
    mem['h049C]=8'h9F; mem['h049D]=8'h04; mem['h049E]=8'h28; mem['h049F]=8'hC5;
    mem['h04A0]=8'hB9; mem['h04A1]=8'h48; mem['h04A2]=8'h98; mem['h04A3]=8'h04;
    mem['h04A4]=8'hC6; mem['h04A5]=8'hBA; mem['h04A6]=8'h48; mem['h04A7]=8'h98;
    mem['h04A8]=8'h04; mem['h04A9]=8'h46; mem['h04AA]=8'h0C; mem['h04AB]=8'h02;
    mem['h04AC]=8'h44; mem['h04AD]=8'hD8; mem['h04AE]=8'h07; mem['h04AF]=8'h46;
    mem['h04B0]=8'h99; mem['h04B1]=8'h02; mem['h04B2]=8'h26; mem['h04B3]=8'h6A;
    mem['h04B4]=8'h46; mem['h04B5]=8'h05; mem['h04B6]=8'h04; mem['h04B7]=8'h46;
    mem['h04B8]=8'h20; mem['h04B9]=8'h03; mem['h04BA]=8'hA0; mem['h04BB]=8'h68;
    mem['h04BC]=8'hC9; mem['h04BD]=8'h04; mem['h04BE]=8'h46; mem['h04BF]=8'h99;
    mem['h04C0]=8'h02; mem['h04C1]=8'h26; mem['h04C2]=8'h6C; mem['h04C3]=8'h46;
    mem['h04C4]=8'h05; mem['h04C5]=8'h04; mem['h04C6]=8'h44; mem['h04C7]=8'hDA;
    mem['h04C8]=8'h04; mem['h04C9]=8'h26; mem['h04CA]=8'h6C; mem['h04CB]=8'h1E;
    mem['h04CC]=8'h6A; mem['h04CD]=8'h46; mem['h04CE]=8'h65; mem['h04CF]=8'h02;
    mem['h04D0]=8'hF4; mem['h04D1]=8'hC7; mem['h04D2]=8'h04; mem['h04D3]=8'hFF;
    mem['h04D4]=8'hF8; mem['h04D5]=8'h30; mem['h04D6]=8'hC7; mem['h04D7]=8'h0C;
    mem['h04D8]=8'h00; mem['h04D9]=8'hF8; mem['h04DA]=8'h1E; mem['h04DB]=8'h6A;
    mem['h04DC]=8'h26; mem['h04DD]=8'h6C; mem['h04DE]=8'h46; mem['h04DF]=8'hE8;
    mem['h04E0]=8'h0D; mem['h04E1]=8'h06; mem['h04E2]=8'h3A; mem['h04E3]=8'h46;
    mem['h04E4]=8'h40; mem['h04E5]=8'h00; mem['h04E6]=8'h06; mem['h04E7]=8'h20;
    mem['h04E8]=8'h46; mem['h04E9]=8'h40; mem['h04EA]=8'h00; mem['h04EB]=8'h46;
    mem['h04EC]=8'h20; mem['h04ED]=8'h03; mem['h04EE]=8'h46; mem['h04EF]=8'hB8;
    mem['h04F0]=8'h02; mem['h04F1]=8'h46; mem['h04F2]=8'hFC; mem['h04F3]=8'h06;
    mem['h04F4]=8'h68; mem['h04F5]=8'hD8; mem['h04F6]=8'h07; mem['h04F7]=8'h46;
    mem['h04F8]=8'h99; mem['h04F9]=8'h02; mem['h04FA]=8'h2E; mem['h04FB]=8'h38;
    mem['h04FC]=8'hF3; mem['h04FD]=8'hC7; mem['h04FE]=8'h24; mem['h04FF]=8'h0F;
    mem['h0500]=8'h48; mem['h0501]=8'hE6; mem['h0502]=8'h04; mem['h0503]=8'h46;
    mem['h0504]=8'h60; mem['h0505]=8'h00; mem['h0506]=8'h44; mem['h0507]=8'hDE;
    mem['h0508]=8'h04; mem['h0509]=8'h2E; mem['h050A]=8'h38; mem['h050B]=8'hF3;
    mem['h050C]=8'h3E; mem['h050D]=8'h00; mem['h050E]=8'h30; mem['h050F]=8'h3E;
    mem['h0510]=8'h00; mem['h0511]=8'h07; mem['h0512]=8'h2E; mem['h0513]=8'h38;
    mem['h0514]=8'hF4; mem['h0515]=8'h3E; mem['h0516]=8'h00; mem['h0517]=8'h30;
    mem['h0518]=8'h3E; mem['h0519]=8'h00; mem['h051A]=8'h07; mem['h051B]=8'h2E;
    mem['h051C]=8'h38; mem['h051D]=8'h3E; mem['h051E]=8'h00; mem['h051F]=8'h30;
    mem['h0520]=8'h3E; mem['h0521]=8'h00; mem['h0522]=8'h07; mem['h0523]=8'h24;
    mem['h0524]=8'h5F; mem['h0525]=8'h14; mem['h0526]=8'h41; mem['h0527]=8'h02;
    mem['h0528]=8'h04; mem['h0529]=8'h02; mem['h052A]=8'h07; mem['h052B]=8'h2E;
    mem['h052C]=8'h38; mem['h052D]=8'hF3; mem['h052E]=8'hF8; mem['h052F]=8'h30;
    mem['h0530]=8'h3E; mem['h0531]=8'h00; mem['h0532]=8'h07; mem['h0533]=8'h2E;
    mem['h0534]=8'h38; mem['h0535]=8'hF3; mem['h0536]=8'hFA; mem['h0537]=8'h30;
    mem['h0538]=8'hF9; mem['h0539]=8'h07; mem['h053A]=8'hF3; mem['h053B]=8'h2E;
    mem['h053C]=8'h38; mem['h053D]=8'hD7; mem['h053E]=8'h30; mem['h053F]=8'hCF;
    mem['h0540]=8'h07; mem['h0541]=8'h2E; mem['h0542]=8'h38; mem['h0543]=8'hF3;
    mem['h0544]=8'h30; mem['h0545]=8'hC7; mem['h0546]=8'h12; mem['h0547]=8'h07;
    mem['h0548]=8'h2E; mem['h0549]=8'h38; mem['h054A]=8'hF3; mem['h054B]=8'hC7;
    mem['h054C]=8'h2C; mem['h054D]=8'hFF; mem['h054E]=8'hF8; mem['h054F]=8'h30;
    mem['h0550]=8'hC7; mem['h0551]=8'h2C; mem['h0552]=8'hFF; mem['h0553]=8'hF8;
    mem['h0554]=8'h44; mem['h0555]=8'h99; mem['h0556]=8'h02; mem['h0557]=8'hF3;
    mem['h0558]=8'h2E; mem['h0559]=8'h38; mem['h055A]=8'hC7; mem['h055B]=8'hA0;
    mem['h055C]=8'h0B; mem['h055D]=8'h30; mem['h055E]=8'hC7; mem['h055F]=8'hA0;
    mem['h0560]=8'h07; mem['h0561]=8'h2E; mem['h0562]=8'h38; mem['h0563]=8'hF0;
    mem['h0564]=8'hC1; mem['h0565]=8'h87; mem['h0566]=8'hF8; mem['h0567]=8'h30;
    mem['h0568]=8'h06; mem['h0569]=8'h00; mem['h056A]=8'h8F; mem['h056B]=8'hF8;
    mem['h056C]=8'h07; mem['h056D]=8'h46; mem['h056E]=8'hCE; mem['h056F]=8'h01;
    mem['h0570]=8'h2E; mem['h0571]=8'h38; mem['h0572]=8'hF4; mem['h0573]=8'hD7;
    mem['h0574]=8'h30; mem['h0575]=8'hCF; mem['h0576]=8'hF3; mem['h0577]=8'hC2;
    mem['h0578]=8'h87; mem['h0579]=8'hF8; mem['h057A]=8'h30; mem['h057B]=8'hC1;
    mem['h057C]=8'h8F; mem['h057D]=8'hF8; mem['h057E]=8'h44; mem['h057F]=8'h0C;
    mem['h0580]=8'h02; mem['h0581]=8'h46; mem['h0582]=8'hCE; mem['h0583]=8'h01;
    mem['h0584]=8'h2E; mem['h0585]=8'h38; mem['h0586]=8'hF3; mem['h0587]=8'hD7;
    mem['h0588]=8'h30; mem['h0589]=8'hCF; mem['h058A]=8'hF4; mem['h058B]=8'hC2;
    mem['h058C]=8'h97; mem['h058D]=8'hD0; mem['h058E]=8'h30; mem['h058F]=8'hC1;
    mem['h0590]=8'h9F; mem['h0591]=8'hC8; mem['h0592]=8'hF3; mem['h0593]=8'hFA;
    mem['h0594]=8'h30; mem['h0595]=8'hF9; mem['h0596]=8'h44; mem['h0597]=8'h0C;
    mem['h0598]=8'h02; mem['h0599]=8'h2E; mem['h059A]=8'h38; mem['h059B]=8'hF0;
    mem['h059C]=8'hA0; mem['h059D]=8'hC7; mem['h059E]=8'h12; mem['h059F]=8'hF8;
    mem['h05A0]=8'h30; mem['h05A1]=8'hC7; mem['h05A2]=8'h12; mem['h05A3]=8'hF8;
    mem['h05A4]=8'h31; mem['h05A5]=8'hC6; mem['h05A6]=8'h07; mem['h05A7]=8'h2E;
    mem['h05A8]=8'h38; mem['h05A9]=8'hF0; mem['h05AA]=8'h30; mem['h05AB]=8'hC7;
    mem['h05AC]=8'hA0; mem['h05AD]=8'h1A; mem['h05AE]=8'hF8; mem['h05AF]=8'h31;
    mem['h05B0]=8'hC7; mem['h05B1]=8'h1A; mem['h05B2]=8'hF8; mem['h05B3]=8'hC6;
    mem['h05B4]=8'h07; mem['h05B5]=8'h46; mem['h05B6]=8'hCE; mem['h05B7]=8'h01;
    mem['h05B8]=8'h46; mem['h05B9]=8'hDE; mem['h05BA]=8'h01; mem['h05BB]=8'h0E;
    mem['h05BC]=8'h56; mem['h05BD]=8'h46; mem['h05BE]=8'h72; mem['h05BF]=8'h02;
    mem['h05C0]=8'h0E; mem['h05C1]=8'h58; mem['h05C2]=8'h46; mem['h05C3]=8'h8C;
    mem['h05C4]=8'h02; mem['h05C5]=8'h2E; mem['h05C6]=8'h38; mem['h05C7]=8'hF3;
    mem['h05C8]=8'h3E; mem['h05C9]=8'h00; mem['h05CA]=8'h30; mem['h05CB]=8'h3E;
    mem['h05CC]=8'h00; mem['h05CD]=8'h26; mem['h05CE]=8'h56; mem['h05CF]=8'h0E;
    mem['h05D0]=8'h58; mem['h05D1]=8'h16; mem['h05D2]=8'h10; mem['h05D3]=8'hC1;
    mem['h05D4]=8'h46; mem['h05D5]=8'hA7; mem['h05D6]=8'h05; mem['h05D7]=8'h40;
    mem['h05D8]=8'hDD; mem['h05D9]=8'h05; mem['h05DA]=8'h46; mem['h05DB]=8'h6D;
    mem['h05DC]=8'h05; mem['h05DD]=8'hC4; mem['h05DE]=8'h46; mem['h05DF]=8'h99;
    mem['h05E0]=8'h05; mem['h05E1]=8'h11; mem['h05E2]=8'h48; mem['h05E3]=8'hD3;
    mem['h05E4]=8'h05; mem['h05E5]=8'h46; mem['h05E6]=8'h1C; mem['h05E7]=8'h02;
    mem['h05E8]=8'h44; mem['h05E9]=8'h0C; mem['h05EA]=8'h02; mem['h05EB]=8'h46;
    mem['h05EC]=8'hCE; mem['h05ED]=8'h01; mem['h05EE]=8'h46; mem['h05EF]=8'hDE;
    mem['h05F0]=8'h01; mem['h05F1]=8'h0E; mem['h05F2]=8'h66; mem['h05F3]=8'h46;
    mem['h05F4]=8'h72; mem['h05F5]=8'h02; mem['h05F6]=8'hD9; mem['h05F7]=8'h0E;
    mem['h05F8]=8'h68; mem['h05F9]=8'h46; mem['h05FA]=8'h8C; mem['h05FB]=8'h02;
    mem['h05FC]=8'hE1; mem['h05FD]=8'h0E; mem['h05FE]=8'h00; mem['h05FF]=8'h16;
    mem['h0600]=8'h01; mem['h0601]=8'h0E; mem['h0602]=8'h00; mem['h0603]=8'h16;
    mem['h0604]=8'h01; mem['h0605]=8'h2E; mem['h0606]=8'h38; mem['h0607]=8'h36;
    mem['h0608]=8'h69; mem['h0609]=8'hC7; mem['h060A]=8'h24; mem['h060B]=8'h80;
    mem['h060C]=8'h48; mem['h060D]=8'h21; mem['h060E]=8'h06; mem['h060F]=8'h06;
    mem['h0610]=8'h68; mem['h0611]=8'h46; mem['h0612]=8'h99; mem['h0613]=8'h05;
    mem['h0614]=8'hA8; mem['h0615]=8'hC2; mem['h0616]=8'h12; mem['h0617]=8'hD0;
    mem['h0618]=8'hC1; mem['h0619]=8'h12; mem['h061A]=8'hC8; mem['h061B]=8'h40;
    mem['h061C]=8'h05; mem['h061D]=8'h06; mem['h061E]=8'h44; mem['h061F]=8'h5F;
    mem['h0620]=8'h06; mem['h0621]=8'h36; mem['h0622]=8'h64; mem['h0623]=8'h46;
    mem['h0624]=8'h1B; mem['h0625]=8'h05; mem['h0626]=8'h1E; mem['h0627]=8'h66;
    mem['h0628]=8'h26; mem['h0629]=8'h68; mem['h062A]=8'h46; mem['h062B]=8'hFC;
    mem['h062C]=8'h06; mem['h062D]=8'h60; mem['h062E]=8'h3E; mem['h062F]=8'h06;
    mem['h0630]=8'h46; mem['h0631]=8'h81; mem['h0632]=8'h05; mem['h0633]=8'h2E;
    mem['h0634]=8'h38; mem['h0635]=8'h36; mem['h0636]=8'h64; mem['h0637]=8'hC2;
    mem['h0638]=8'h87; mem['h0639]=8'hF8; mem['h063A]=8'h30; mem['h063B]=8'hC1;
    mem['h063C]=8'h8F; mem['h063D]=8'hF8; mem['h063E]=8'h06; mem['h063F]=8'h68;
    mem['h0640]=8'h46; mem['h0641]=8'hA7; mem['h0642]=8'h05; mem['h0643]=8'hA8;
    mem['h0644]=8'hC1; mem['h0645]=8'h1A; mem['h0646]=8'hC8; mem['h0647]=8'hC2;
    mem['h0648]=8'h1A; mem['h0649]=8'hD0; mem['h064A]=8'h40; mem['h064B]=8'h26;
    mem['h064C]=8'h06; mem['h064D]=8'h1E; mem['h064E]=8'h46; mem['h064F]=8'h26;
    mem['h0650]=8'h66; mem['h0651]=8'h46; mem['h0652]=8'h58; mem['h0653]=8'h02;
    mem['h0654]=8'h46; mem['h0655]=8'h1C; mem['h0656]=8'h02; mem['h0657]=8'h0E;
    mem['h0658]=8'h64; mem['h0659]=8'h46; mem['h065A]=8'h7F; mem['h065B]=8'h02;
    mem['h065C]=8'h44; mem['h065D]=8'h0C; mem['h065E]=8'h02; mem['h065F]=8'h2E;
    mem['h0660]=8'h38; mem['h0661]=8'h36; mem['h0662]=8'h46; mem['h0663]=8'h3E;
    mem['h0664]=8'h00; mem['h0665]=8'h30; mem['h0666]=8'h3E; mem['h0667]=8'h00;
    mem['h0668]=8'h36; mem['h0669]=8'h64; mem['h066A]=8'h3E; mem['h066B]=8'hFF;
    mem['h066C]=8'h30; mem['h066D]=8'h3E; mem['h066E]=8'h7F; mem['h066F]=8'h44;
    mem['h0670]=8'h54; mem['h0671]=8'h06; mem['h0672]=8'hC4; mem['h0673]=8'h46;
    mem['h0674]=8'h2C; mem['h0675]=8'h02; mem['h0676]=8'h46; mem['h0677]=8'hCE;
    mem['h0678]=8'h01; mem['h0679]=8'hD3; mem['h067A]=8'h2E; mem['h067B]=8'h38;
    mem['h067C]=8'h36; mem['h067D]=8'h71; mem['h067E]=8'h3E; mem['h067F]=8'h00;
    mem['h0680]=8'h2E; mem['h0681]=8'h38; mem['h0682]=8'h36; mem['h0683]=8'h72;
    mem['h0684]=8'h3E; mem['h0685]=8'h00; mem['h0686]=8'h46; mem['h0687]=8'h41;
    mem['h0688]=8'h05; mem['h0689]=8'h40; mem['h068A]=8'h95; mem['h068B]=8'h06;
    mem['h068C]=8'h46; mem['h068D]=8'h48; mem['h068E]=8'h05; mem['h068F]=8'h2E;
    mem['h0690]=8'h38; mem['h0691]=8'h36; mem['h0692]=8'h71; mem['h0693]=8'h3E;
    mem['h0694]=8'h01; mem['h0695]=8'hDC; mem['h0696]=8'h46; mem['h0697]=8'h41;
    mem['h0698]=8'h05; mem['h0699]=8'h40; mem['h069A]=8'hA5; mem['h069B]=8'h06;
    mem['h069C]=8'h46; mem['h069D]=8'h48; mem['h069E]=8'h05; mem['h069F]=8'h2E;
    mem['h06A0]=8'h38; mem['h06A1]=8'h36; mem['h06A2]=8'h72; mem['h06A3]=8'h3E;
    mem['h06A4]=8'h01; mem['h06A5]=8'hDA; mem['h06A6]=8'h46; mem['h06A7]=8'hEB;
    mem['h06A8]=8'h05; mem['h06A9]=8'h2E; mem['h06AA]=8'h38; mem['h06AB]=8'h36;
    mem['h06AC]=8'h71; mem['h06AD]=8'hC7; mem['h06AE]=8'hA0; mem['h06AF]=8'h68;
    mem['h06B0]=8'hB7; mem['h06B1]=8'h06; mem['h06B2]=8'h1E; mem['h06B3]=8'h46;
    mem['h06B4]=8'h46; mem['h06B5]=8'h48; mem['h06B6]=8'h05; mem['h06B7]=8'h2E;
    mem['h06B8]=8'h38; mem['h06B9]=8'h36; mem['h06BA]=8'h71; mem['h06BB]=8'hC7;
    mem['h06BC]=8'h2E; mem['h06BD]=8'h38; mem['h06BE]=8'h36; mem['h06BF]=8'h72;
    mem['h06C0]=8'hBF; mem['h06C1]=8'h68; mem['h06C2]=8'hC8; mem['h06C3]=8'h06;
    mem['h06C4]=8'hDA; mem['h06C5]=8'h46; mem['h06C6]=8'h48; mem['h06C7]=8'h05;
    mem['h06C8]=8'h46; mem['h06C9]=8'h0C; mem['h06CA]=8'h02; mem['h06CB]=8'hC4;
    mem['h06CC]=8'h44; mem['h06CD]=8'h42; mem['h06CE]=8'h02; mem['h06CF]=8'h2E;
    mem['h06D0]=8'h38; mem['h06D1]=8'hF4; mem['h06D2]=8'hC7; mem['h06D3]=8'hF3;
    mem['h06D4]=8'hAF; mem['h06D5]=8'hF8; mem['h06D6]=8'hF4; mem['h06D7]=8'h30;
    mem['h06D8]=8'hC7; mem['h06D9]=8'hF3; mem['h06DA]=8'h30; mem['h06DB]=8'hAF;
    mem['h06DC]=8'hF8; mem['h06DD]=8'h07; mem['h06DE]=8'h2E; mem['h06DF]=8'h38;
    mem['h06E0]=8'hF4; mem['h06E1]=8'hC7; mem['h06E2]=8'hF3; mem['h06E3]=8'hA7;
    mem['h06E4]=8'hF8; mem['h06E5]=8'hF4; mem['h06E6]=8'h30; mem['h06E7]=8'hC7;
    mem['h06E8]=8'hF3; mem['h06E9]=8'h30; mem['h06EA]=8'hA7; mem['h06EB]=8'hF8;
    mem['h06EC]=8'h07; mem['h06ED]=8'h2E; mem['h06EE]=8'h38; mem['h06EF]=8'hF4;
    mem['h06F0]=8'hC7; mem['h06F1]=8'hF3; mem['h06F2]=8'hB7; mem['h06F3]=8'hF8;
    mem['h06F4]=8'hF4; mem['h06F5]=8'h30; mem['h06F6]=8'hC7; mem['h06F7]=8'hF3;
    mem['h06F8]=8'h30; mem['h06F9]=8'hB7; mem['h06FA]=8'hF8; mem['h06FB]=8'h07;
    mem['h06FC]=8'h2E; mem['h06FD]=8'h38; mem['h06FE]=8'hF3; mem['h06FF]=8'h30;
    mem['h0700]=8'hC7; mem['h0701]=8'hF4; mem['h0702]=8'h30; mem['h0703]=8'hBF;
    mem['h0704]=8'h0B; mem['h0705]=8'hF3; mem['h0706]=8'hC7; mem['h0707]=8'hF4;
    mem['h0708]=8'hBF; mem['h0709]=8'h07; mem['h070A]=8'h2E; mem['h070B]=8'h38;
    mem['h070C]=8'hF3; mem['h070D]=8'h30; mem['h070E]=8'hC7; mem['h070F]=8'h12;
    mem['h0710]=8'h60; mem['h0711]=8'h1D; mem['h0712]=8'h07; mem['h0713]=8'hF4;
    mem['h0714]=8'h30; mem['h0715]=8'hC7; mem['h0716]=8'h12; mem['h0717]=8'h60;
    mem['h0718]=8'h2F; mem['h0719]=8'h07; mem['h071A]=8'h44; mem['h071B]=8'hFC;
    mem['h071C]=8'h06; mem['h071D]=8'hF4; mem['h071E]=8'h30; mem['h071F]=8'hC7;
    mem['h0720]=8'h12; mem['h0721]=8'h40; mem['h0722]=8'h33; mem['h0723]=8'h07;
    mem['h0724]=8'h46; mem['h0725]=8'hFC; mem['h0726]=8'h06; mem['h0727]=8'h2B;
    mem['h0728]=8'h06; mem['h0729]=8'h01; mem['h072A]=8'h12; mem['h072B]=8'h2C;
    mem['h072C]=8'h01; mem['h072D]=8'h1A; mem['h072E]=8'h07; mem['h072F]=8'hA8;
    mem['h0730]=8'h04; mem['h0731]=8'h01; mem['h0732]=8'h07; mem['h0733]=8'hA8;
    mem['h0734]=8'h14; mem['h0735]=8'h01; mem['h0736]=8'h07; mem['h0737]=8'h46;
    mem['h0738]=8'hCE; mem['h0739]=8'h01; mem['h073A]=8'h46; mem['h073B]=8'hDE;
    mem['h073C]=8'h01; mem['h073D]=8'h1E; mem['h073E]=8'h52; mem['h073F]=8'h26;
    mem['h0740]=8'h4A; mem['h0741]=8'h46; mem['h0742]=8'h58; mem['h0743]=8'h02;
    mem['h0744]=8'hC3; mem['h0745]=8'h46; mem['h0746]=8'h99; mem['h0747]=8'h05;
    mem['h0748]=8'h46; mem['h0749]=8'h99; mem['h074A]=8'h05; mem['h074B]=8'h46;
    mem['h074C]=8'h99; mem['h074D]=8'h05; mem['h074E]=8'h46; mem['h074F]=8'h99;
    mem['h0750]=8'h05; mem['h0751]=8'h46; mem['h0752]=8'h99; mem['h0753]=8'h05;
    mem['h0754]=8'h46; mem['h0755]=8'hCF; mem['h0756]=8'h06; mem['h0757]=8'h1E;
    mem['h0758]=8'h4C; mem['h0759]=8'h46; mem['h075A]=8'h65; mem['h075B]=8'h02;
    mem['h075C]=8'h1E; mem['h075D]=8'h54; mem['h075E]=8'h26; mem['h075F]=8'h52;
    mem['h0760]=8'h46; mem['h0761]=8'h58; mem['h0762]=8'h02; mem['h0763]=8'hC3;
    mem['h0764]=8'h46; mem['h0765]=8'hA7; mem['h0766]=8'h05; mem['h0767]=8'h46;
    mem['h0768]=8'hA7; mem['h0769]=8'h05; mem['h076A]=8'h46; mem['h076B]=8'hA7;
    mem['h076C]=8'h05; mem['h076D]=8'h46; mem['h076E]=8'hCF; mem['h076F]=8'h06;
    mem['h0770]=8'h1E; mem['h0771]=8'h4C; mem['h0772]=8'h26; mem['h0773]=8'h52;
    mem['h0774]=8'h46; mem['h0775]=8'h65; mem['h0776]=8'h02; mem['h0777]=8'hC4;
    mem['h0778]=8'h46; mem['h0779]=8'hA7; mem['h077A]=8'h05; mem['h077B]=8'h46;
    mem['h077C]=8'hCF; mem['h077D]=8'h06; mem['h077E]=8'h26; mem['h077F]=8'h54;
    mem['h0780]=8'h46; mem['h0781]=8'hCF; mem['h0782]=8'h06; mem['h0783]=8'h46;
    mem['h0784]=8'h1C; mem['h0785]=8'h02; mem['h0786]=8'h44; mem['h0787]=8'h0C;
    mem['h0788]=8'h02; mem['h0789]=8'h2E; mem['h078A]=8'h3F; mem['h078B]=8'h36;
    mem['h078C]=8'h00; mem['h078D]=8'h3E; mem['h078E]=8'h00; mem['h078F]=8'h2E;
    mem['h0790]=8'h3E; mem['h0791]=8'h36; mem['h0792]=8'h00; mem['h0793]=8'h3E;
    mem['h0794]=8'h00; mem['h0795]=8'h2E; mem['h0796]=8'h38; mem['h0797]=8'h36;
    mem['h0798]=8'h74; mem['h0799]=8'h3E; mem['h079A]=8'h10; mem['h079B]=8'h30;
    mem['h079C]=8'h3E; mem['h079D]=8'h27; mem['h079E]=8'h30; mem['h079F]=8'h3E;
    mem['h07A0]=8'hE8; mem['h07A1]=8'h30; mem['h07A2]=8'h3E; mem['h07A3]=8'h03;
    mem['h07A4]=8'h30; mem['h07A5]=8'h3E; mem['h07A6]=8'h64; mem['h07A7]=8'h30;
    mem['h07A8]=8'h3E; mem['h07A9]=8'h00; mem['h07AA]=8'h30; mem['h07AB]=8'h3E;
    mem['h07AC]=8'h0A; mem['h07AD]=8'h30; mem['h07AE]=8'h3E; mem['h07AF]=8'h00;
    mem['h07B0]=8'h2E; mem['h07B1]=8'h01; mem['h07B2]=8'h36; mem['h07B3]=8'h0F;
    mem['h07B4]=8'h46; mem['h07B5]=8'h52; mem['h07B6]=8'h00; mem['h07B7]=8'h2E;
    mem['h07B8]=8'h38; mem['h07B9]=8'h36; mem['h07BA]=8'h3C; mem['h07BB]=8'h3E;
    mem['h07BC]=8'h00; mem['h07BD]=8'h30; mem['h07BE]=8'h3E; mem['h07BF]=8'h10;
    mem['h07C0]=8'h31; mem['h07C1]=8'h2E; mem['h07C2]=8'h38; mem['h07C3]=8'h36;
    mem['h07C4]=8'h4A; mem['h07C5]=8'h3E; mem['h07C6]=8'hD2; mem['h07C7]=8'h30;
    mem['h07C8]=8'h3E; mem['h07C9]=8'h04; mem['h07CA]=8'h31; mem['h07CB]=8'h2E;
    mem['h07CC]=8'h38; mem['h07CD]=8'h36; mem['h07CE]=8'h4C; mem['h07CF]=8'h3E;
    mem['h07D0]=8'hD2; mem['h07D1]=8'h30; mem['h07D2]=8'h3E; mem['h07D3]=8'h04;
    mem['h07D4]=8'h31; mem['h07D5]=8'h44; mem['h07D6]=8'h22; mem['h07D7]=8'h08;
    mem['h07D8]=8'h2E; mem['h07D9]=8'h38; mem['h07DA]=8'h36; mem['h07DB]=8'h6E;
    mem['h07DC]=8'h46; mem['h07DD]=8'h58; mem['h07DE]=8'h05; mem['h07DF]=8'h68;
    mem['h07E0]=8'h22; mem['h07E1]=8'h08; mem['h07E2]=8'h1E; mem['h07E3]=8'h6E;
    mem['h07E4]=8'h46; mem['h07E5]=8'h94; mem['h07E6]=8'h0E; mem['h07E7]=8'h06;
    mem['h07E8]=8'h20; mem['h07E9]=8'h46; mem['h07EA]=8'h40; mem['h07EB]=8'h00;
    mem['h07EC]=8'h2E; mem['h07ED]=8'h38; mem['h07EE]=8'h36; mem['h07EF]=8'h70;
    mem['h07F0]=8'hC7; mem['h07F1]=8'h46; mem['h07F2]=8'hB8; mem['h07F3]=8'h02;
    mem['h07F4]=8'h06; mem['h07F5]=8'h20; mem['h07F6]=8'h46; mem['h07F7]=8'h40;
    mem['h07F8]=8'h00; mem['h07F9]=8'h2E; mem['h07FA]=8'h01; mem['h07FB]=8'h36;
    mem['h07FC]=8'h6A; mem['h07FD]=8'h46; mem['h07FE]=8'h52; mem['h07FF]=8'h00;
    mem['h0800]=8'h1E; mem['h0801]=8'h00; mem['h0802]=8'h46; mem['h0803]=8'hA5;
    mem['h0804]=8'h02; mem['h0805]=8'h46; mem['h0806]=8'h94; mem['h0807]=8'h0E;
    mem['h0808]=8'h46; mem['h0809]=8'h60; mem['h080A]=8'h00; mem['h080B]=8'h1E;
    mem['h080C]=8'h36; mem['h080D]=8'h46; mem['h080E]=8'h57; mem['h080F]=8'h05;
    mem['h0810]=8'h68; mem['h0811]=8'h22; mem['h0812]=8'h08; mem['h0813]=8'h2E;
    mem['h0814]=8'h01; mem['h0815]=8'h36; mem['h0816]=8'h79; mem['h0817]=8'h46;
    mem['h0818]=8'h52; mem['h0819]=8'h00; mem['h081A]=8'h1E; mem['h081B]=8'h36;
    mem['h081C]=8'h46; mem['h081D]=8'h66; mem['h081E]=8'h0D; mem['h081F]=8'h46;
    mem['h0820]=8'h60; mem['h0821]=8'h00; mem['h0822]=8'h2E; mem['h0823]=8'h3F;
    mem['h0824]=8'h36; mem['h0825]=8'h00; mem['h0826]=8'hC7; mem['h0827]=8'hD0;
    mem['h0828]=8'hA0; mem['h0829]=8'h68; mem['h082A]=8'h3A; mem['h082B]=8'h08;
    mem['h082C]=8'h2E; mem['h082D]=8'h01; mem['h082E]=8'h36; mem['h082F]=8'h6F;
    mem['h0830]=8'h46; mem['h0831]=8'h52; mem['h0832]=8'h00; mem['h0833]=8'hC2;
    mem['h0834]=8'h46; mem['h0835]=8'hB8; mem['h0836]=8'h02; mem['h0837]=8'h46;
    mem['h0838]=8'h60; mem['h0839]=8'h00; mem['h083A]=8'h2E; mem['h083B]=8'h3E;
    mem['h083C]=8'h36; mem['h083D]=8'h00; mem['h083E]=8'hC7; mem['h083F]=8'hD0;
    mem['h0840]=8'hA0; mem['h0841]=8'h68; mem['h0842]=8'h52; mem['h0843]=8'h08;
    mem['h0844]=8'h2E; mem['h0845]=8'h01; mem['h0846]=8'h36; mem['h0847]=8'h73;
    mem['h0848]=8'h46; mem['h0849]=8'h52; mem['h084A]=8'h00; mem['h084B]=8'hC2;
    mem['h084C]=8'h46; mem['h084D]=8'hB8; mem['h084E]=8'h02; mem['h084F]=8'h46;
    mem['h0850]=8'h60; mem['h0851]=8'h00; mem['h0852]=8'hA8; mem['h0853]=8'h2E;
    mem['h0854]=8'h3F; mem['h0855]=8'h36; mem['h0856]=8'h00; mem['h0857]=8'hF8;
    mem['h0858]=8'h2E; mem['h0859]=8'h3E; mem['h085A]=8'h36; mem['h085B]=8'h00;
    mem['h085C]=8'hF8; mem['h085D]=8'h2E; mem['h085E]=8'h38; mem['h085F]=8'h36;
    mem['h0860]=8'h48; mem['h0861]=8'h3E; mem['h0862]=8'h00; mem['h0863]=8'h30;
    mem['h0864]=8'h3E; mem['h0865]=8'h3D; mem['h0866]=8'h31; mem['h0867]=8'hA8;
    mem['h0868]=8'h2E; mem['h0869]=8'h38; mem['h086A]=8'h36; mem['h086B]=8'h6E;
    mem['h086C]=8'hF8; mem['h086D]=8'h30; mem['h086E]=8'hF8; mem['h086F]=8'h36;
    mem['h0870]=8'h70; mem['h0871]=8'hF8; mem['h0872]=8'h2E; mem['h0873]=8'h01;
    mem['h0874]=8'h36; mem['h0875]=8'h44; mem['h0876]=8'h46; mem['h0877]=8'h52;
    mem['h0878]=8'h00; mem['h0879]=8'h36; mem['h087A]=8'h36; mem['h087B]=8'h46;
    mem['h087C]=8'h1B; mem['h087D]=8'h05; mem['h087E]=8'h2E; mem['h087F]=8'h38;
    mem['h0880]=8'h36; mem['h0881]=8'h00; mem['h0882]=8'h3E; mem['h0883]=8'h00;
    mem['h0884]=8'h30; mem['h0885]=8'h3E; mem['h0886]=8'h3D; mem['h0887]=8'h31;
    mem['h0888]=8'h1E; mem['h0889]=8'h00; mem['h088A]=8'h46; mem['h088B]=8'hA8;
    mem['h088C]=8'h03; mem['h088D]=8'h46; mem['h088E]=8'h20; mem['h088F]=8'h03;
    mem['h0890]=8'h3C; mem['h0891]=8'h2E; mem['h0892]=8'h68; mem['h0893]=8'h7A;
    mem['h0894]=8'h04; mem['h0895]=8'h46; mem['h0896]=8'hE0; mem['h0897]=8'h02;
    mem['h0898]=8'h60; mem['h0899]=8'hD0; mem['h089A]=8'h0C; mem['h089B]=8'h2E;
    mem['h089C]=8'h38; mem['h089D]=8'h36; mem['h089E]=8'h36; mem['h089F]=8'h3E;
    mem['h08A0]=8'h00; mem['h08A1]=8'h30; mem['h08A2]=8'h3E; mem['h08A3]=8'h00;
    mem['h08A4]=8'h31; mem['h08A5]=8'h2E; mem['h08A6]=8'h38; mem['h08A7]=8'h36;
    mem['h08A8]=8'h3A; mem['h08A9]=8'h3E; mem['h08AA]=8'hFF; mem['h08AB]=8'h30;
    mem['h08AC]=8'h3E; mem['h08AD]=8'h37; mem['h08AE]=8'h31; mem['h08AF]=8'h1E;
    mem['h08B0]=8'h00; mem['h08B1]=8'h44; mem['h08B2]=8'h4A; mem['h08B3]=8'h09;
    mem['h08B4]=8'h2E; mem['h08B5]=8'h38; mem['h08B6]=8'h36; mem['h08B7]=8'h00;
    mem['h08B8]=8'h3E; mem['h08B9]=8'h00; mem['h08BA]=8'h30; mem['h08BB]=8'h3E;
    mem['h08BC]=8'h10; mem['h08BD]=8'h31; mem['h08BE]=8'hDE; mem['h08BF]=8'h26;
    mem['h08C0]=8'h38; mem['h08C1]=8'h46; mem['h08C2]=8'h65; mem['h08C3]=8'h02;
    mem['h08C4]=8'h26; mem['h08C5]=8'h52; mem['h08C6]=8'h46; mem['h08C7]=8'h68;
    mem['h08C8]=8'h03; mem['h08C9]=8'h46; mem['h08CA]=8'h99; mem['h08CB]=8'h02;
    mem['h08CC]=8'h46; mem['h08CD]=8'h99; mem['h08CE]=8'h02; mem['h08CF]=8'h1E;
    mem['h08D0]=8'h52; mem['h08D1]=8'h26; mem['h08D2]=8'h36; mem['h08D3]=8'h46;
    mem['h08D4]=8'hFC; mem['h08D5]=8'h06; mem['h08D6]=8'h40; mem['h08D7]=8'hEB;
    mem['h08D8]=8'h08; mem['h08D9]=8'h1E; mem['h08DA]=8'h00; mem['h08DB]=8'h26;
    mem['h08DC]=8'h00; mem['h08DD]=8'h46; mem['h08DE]=8'h68; mem['h08DF]=8'h03;
    mem['h08E0]=8'h26; mem['h08E1]=8'h3C; mem['h08E2]=8'h46; mem['h08E3]=8'hFC;
    mem['h08E4]=8'h06; mem['h08E5]=8'h60; mem['h08E6]=8'hBF; mem['h08E7]=8'h08;
    mem['h08E8]=8'h44; mem['h08E9]=8'hD8; mem['h08EA]=8'h07; mem['h08EB]=8'h46;
    mem['h08EC]=8'h65; mem['h08ED]=8'h02; mem['h08EE]=8'h44; mem['h08EF]=8'h03;
    mem['h08F0]=8'h09; mem['h08F1]=8'h1E; mem['h08F2]=8'h00; mem['h08F3]=8'h26;
    mem['h08F4]=8'h38; mem['h08F5]=8'h46; mem['h08F6]=8'h65; mem['h08F7]=8'h02;
    mem['h08F8]=8'h26; mem['h08F9]=8'h36; mem['h08FA]=8'h46; mem['h08FB]=8'h68;
    mem['h08FC]=8'h03; mem['h08FD]=8'h46; mem['h08FE]=8'h99; mem['h08FF]=8'h02;
    mem['h0900]=8'h46; mem['h0901]=8'h99; mem['h0902]=8'h02; mem['h0903]=8'h1E;
    mem['h0904]=8'h00; mem['h0905]=8'h26; mem['h0906]=8'h3A; mem['h0907]=8'h46;
    mem['h0908]=8'h68; mem['h0909]=8'h03; mem['h090A]=8'h46; mem['h090B]=8'h99;
    mem['h090C]=8'h02; mem['h090D]=8'h46; mem['h090E]=8'h99; mem['h090F]=8'h02;
    mem['h0910]=8'h44; mem['h0911]=8'h4A; mem['h0912]=8'h09; mem['h0913]=8'h1E;
    mem['h0914]=8'h48; mem['h0915]=8'h26; mem['h0916]=8'h3A; mem['h0917]=8'h46;
    mem['h0918]=8'h68; mem['h0919]=8'h03; mem['h091A]=8'h46; mem['h091B]=8'h99;
    mem['h091C]=8'h02; mem['h091D]=8'h46; mem['h091E]=8'h99; mem['h091F]=8'h02;
    mem['h0920]=8'h26; mem['h0921]=8'h38; mem['h0922]=8'h46; mem['h0923]=8'h68;
    mem['h0924]=8'h03; mem['h0925]=8'h46; mem['h0926]=8'h99; mem['h0927]=8'h02;
    mem['h0928]=8'h46; mem['h0929]=8'h99; mem['h092A]=8'h02; mem['h092B]=8'h26;
    mem['h092C]=8'h00; mem['h092D]=8'h46; mem['h092E]=8'h68; mem['h092F]=8'h03;
    mem['h0930]=8'h46; mem['h0931]=8'h99; mem['h0932]=8'h02; mem['h0933]=8'h46;
    mem['h0934]=8'h99; mem['h0935]=8'h02; mem['h0936]=8'h1E; mem['h0937]=8'h3A;
    mem['h0938]=8'h26; mem['h0939]=8'h3C; mem['h093A]=8'h46; mem['h093B]=8'hFC;
    mem['h093C]=8'h06; mem['h093D]=8'h40; mem['h093E]=8'hD8; mem['h093F]=8'h07;
    mem['h0940]=8'h1E; mem['h0941]=8'h00; mem['h0942]=8'h26; mem['h0943]=8'h3A;
    mem['h0944]=8'h46; mem['h0945]=8'h58; mem['h0946]=8'h02; mem['h0947]=8'h44;
    mem['h0948]=8'hF1; mem['h0949]=8'h08; mem['h094A]=8'h1E; mem['h094B]=8'h00;
    mem['h094C]=8'h46; mem['h094D]=8'h20; mem['h094E]=8'h03; mem['h094F]=8'h3C;
    mem['h0950]=8'h20; mem['h0951]=8'h48; mem['h0952]=8'h5A; mem['h0953]=8'h09;
    mem['h0954]=8'h46; mem['h0955]=8'h99; mem['h0956]=8'h02; mem['h0957]=8'h44;
    mem['h0958]=8'h4C; mem['h0959]=8'h09; mem['h095A]=8'hA0; mem['h095B]=8'h68;
    mem['h095C]=8'h36; mem['h095D]=8'h09; mem['h095E]=8'h46; mem['h095F]=8'h99;
    mem['h0960]=8'h02; mem['h0961]=8'h3C; mem['h0962]=8'h3F; mem['h0963]=8'h68;
    mem['h0964]=8'hDD; mem['h0965]=8'h09; mem['h0966]=8'h3C; mem['h0967]=8'h5D;
    mem['h0968]=8'h68; mem['h0969]=8'h13; mem['h096A]=8'h09; mem['h096B]=8'h3C;
    mem['h096C]=8'h40; mem['h096D]=8'h48; mem['h096E]=8'h7D; mem['h096F]=8'h09;
    mem['h0970]=8'h0E; mem['h0971]=8'h09; mem['h0972]=8'h16; mem['h0973]=8'h79;
    mem['h0974]=8'h26; mem['h0975]=8'h4E; mem['h0976]=8'h44; mem['h0977]=8'hA9;
    mem['h0978]=8'h0B; mem['h0979]=8'h1E; mem['h097A]=8'h00; mem['h097B]=8'h06;
    mem['h097C]=8'h40; mem['h097D]=8'h46; mem['h097E]=8'hB0; mem['h097F]=8'h01;
    mem['h0980]=8'h46; mem['h0981]=8'h20; mem['h0982]=8'h03; mem['h0983]=8'h3C;
    mem['h0984]=8'h3D; mem['h0985]=8'h68; mem['h0986]=8'h8E; mem['h0987]=8'h09;
    mem['h0988]=8'h46; mem['h0989]=8'hEE; mem['h098A]=8'h01; mem['h098B]=8'h44;
    mem['h098C]=8'hCB; mem['h098D]=8'h09; mem['h098E]=8'h46; mem['h098F]=8'h99;
    mem['h0990]=8'h02; mem['h0991]=8'h0E; mem['h0992]=8'h09; mem['h0993]=8'h16;
    mem['h0994]=8'h9A; mem['h0995]=8'h26; mem['h0996]=8'h44; mem['h0997]=8'h44;
    mem['h0998]=8'h87; mem['h0999]=8'h0A; mem['h099A]=8'h46; mem['h099B]=8'hEE;
    mem['h099C]=8'h01; mem['h099D]=8'h46; mem['h099E]=8'h04; mem['h099F]=8'h03;
    mem['h09A0]=8'h60; mem['h09A1]=8'hED; mem['h09A2]=8'h09; mem['h09A3]=8'h3C;
    mem['h09A4]=8'h40; mem['h09A5]=8'h68; mem['h09A6]=8'hF9; mem['h09A7]=8'h09;
    mem['h09A8]=8'h3C; mem['h09A9]=8'h3B; mem['h09AA]=8'h68; mem['h09AB]=8'h16;
    mem['h09AC]=8'h0A; mem['h09AD]=8'h3C; mem['h09AE]=8'h23; mem['h09AF]=8'h68;
    mem['h09B0]=8'h21; mem['h09B1]=8'h0A; mem['h09B2]=8'h3C; mem['h09B3]=8'h21;
    mem['h09B4]=8'h68; mem['h09B5]=8'h61; mem['h09B6]=8'h0A; mem['h09B7]=8'h3C;
    mem['h09B8]=8'h26; mem['h09B9]=8'h68; mem['h09BA]=8'h33; mem['h09BB]=8'h0A;
    mem['h09BC]=8'h3C; mem['h09BD]=8'h24; mem['h09BE]=8'h68; mem['h09BF]=8'h3D;
    mem['h09C0]=8'h0A; mem['h09C1]=8'h3C; mem['h09C2]=8'h27; mem['h09C3]=8'h68;
    mem['h09C4]=8'h48; mem['h09C5]=8'h0A; mem['h09C6]=8'h3C; mem['h09C7]=8'h3E;
    mem['h09C8]=8'h68; mem['h09C9]=8'h57; mem['h09CA]=8'h0A; mem['h09CB]=8'h2E;
    mem['h09CC]=8'h38; mem['h09CD]=8'h36; mem['h09CE]=8'h70; mem['h09CF]=8'hF8;
    mem['h09D0]=8'h2E; mem['h09D1]=8'h38; mem['h09D2]=8'h36; mem['h09D3]=8'h6E;
    mem['h09D4]=8'h3E; mem['h09D5]=8'h4B; mem['h09D6]=8'h30; mem['h09D7]=8'h3E;
    mem['h09D8]=8'h01; mem['h09D9]=8'h31; mem['h09DA]=8'h44; mem['h09DB]=8'hD8;
    mem['h09DC]=8'h07; mem['h09DD]=8'h46; mem['h09DE]=8'h20; mem['h09DF]=8'h03;
    mem['h09E0]=8'h3C; mem['h09E1]=8'h24; mem['h09E2]=8'h68; mem['h09E3]=8'h55;
    mem['h09E4]=8'h0E; mem['h09E5]=8'h3C; mem['h09E6]=8'h3F; mem['h09E7]=8'h68;
    mem['h09E8]=8'h77; mem['h09E9]=8'h0E; mem['h09EA]=8'h44; mem['h09EB]=8'h06;
    mem['h09EC]=8'h0E; mem['h09ED]=8'h46; mem['h09EE]=8'h23; mem['h09EF]=8'h05;
    mem['h09F0]=8'hE0; mem['h09F1]=8'h1E; mem['h09F2]=8'h44; mem['h09F3]=8'h46;
    mem['h09F4]=8'h65; mem['h09F5]=8'h02; mem['h09F6]=8'h44; mem['h09F7]=8'h4A;
    mem['h09F8]=8'h09; mem['h09F9]=8'h1E; mem['h09FA]=8'h4E; mem['h09FB]=8'hC3;
    mem['h09FC]=8'h46; mem['h09FD]=8'h99; mem['h09FE]=8'h05; mem['h09FF]=8'h26;
    mem['h0A00]=8'h52; mem['h0A01]=8'h2E; mem['h0A02]=8'h38; mem['h0A03]=8'hF4;
    mem['h0A04]=8'h3E; mem['h0A05]=8'h00; mem['h0A06]=8'h30; mem['h0A07]=8'h3E;
    mem['h0A08]=8'h39; mem['h0A09]=8'h46; mem['h0A0A]=8'h6D; mem['h0A0B]=8'h05;
    mem['h0A0C]=8'h1E; mem['h0A0D]=8'h4E; mem['h0A0E]=8'h26; mem['h0A0F]=8'h44;
    mem['h0A10]=8'h46; mem['h0A11]=8'h89; mem['h0A12]=8'h03; mem['h0A13]=8'h44;
    mem['h0A14]=8'h4A; mem['h0A15]=8'h09; mem['h0A16]=8'h1E; mem['h0A17]=8'h44;
    mem['h0A18]=8'h46; mem['h0A19]=8'h57; mem['h0A1A]=8'h05; mem['h0A1B]=8'h68;
    mem['h0A1C]=8'h36; mem['h0A1D]=8'h09; mem['h0A1E]=8'h44; mem['h0A1F]=8'h4A;
    mem['h0A20]=8'h09; mem['h0A21]=8'h1E; mem['h0A22]=8'h44; mem['h0A23]=8'h46;
    mem['h0A24]=8'h57; mem['h0A25]=8'h05; mem['h0A26]=8'h68; mem['h0A27]=8'h4A;
    mem['h0A28]=8'h09; mem['h0A29]=8'h1E; mem['h0A2A]=8'h36; mem['h0A2B]=8'h26;
    mem['h0A2C]=8'h44; mem['h0A2D]=8'h46; mem['h0A2E]=8'h58; mem['h0A2F]=8'h02;
    mem['h0A30]=8'h44; mem['h0A31]=8'hB4; mem['h0A32]=8'h08; mem['h0A33]=8'h1E;
    mem['h0A34]=8'h3C; mem['h0A35]=8'h26; mem['h0A36]=8'h44; mem['h0A37]=8'h46;
    mem['h0A38]=8'h58; mem['h0A39]=8'h02; mem['h0A3A]=8'h44; mem['h0A3B]=8'h4A;
    mem['h0A3C]=8'h09; mem['h0A3D]=8'h2E; mem['h0A3E]=8'h38; mem['h0A3F]=8'h36;
    mem['h0A40]=8'h44; mem['h0A41]=8'hC7; mem['h0A42]=8'h46; mem['h0A43]=8'h40;
    mem['h0A44]=8'h00; mem['h0A45]=8'h44; mem['h0A46]=8'h4A; mem['h0A47]=8'h09;
    mem['h0A48]=8'h26; mem['h0A49]=8'h44; mem['h0A4A]=8'h1E; mem['h0A4B]=8'h4A;
    mem['h0A4C]=8'h46; mem['h0A4D]=8'h58; mem['h0A4E]=8'h02; mem['h0A4F]=8'h1E;
    mem['h0A50]=8'h4C; mem['h0A51]=8'h46; mem['h0A52]=8'h58; mem['h0A53]=8'h02;
    mem['h0A54]=8'h44; mem['h0A55]=8'h4A; mem['h0A56]=8'h09; mem['h0A57]=8'h26;
    mem['h0A58]=8'h44; mem['h0A59]=8'h1E; mem['h0A5A]=8'h00; mem['h0A5B]=8'h46;
    mem['h0A5C]=8'h58; mem['h0A5D]=8'h02; mem['h0A5E]=8'h44; mem['h0A5F]=8'hF1;
    mem['h0A60]=8'h08; mem['h0A61]=8'h1E; mem['h0A62]=8'h48; mem['h0A63]=8'h26;
    mem['h0A64]=8'h00; mem['h0A65]=8'h46; mem['h0A66]=8'hA5; mem['h0A67]=8'h02;
    mem['h0A68]=8'h46; mem['h0A69]=8'hA5; mem['h0A6A]=8'h02; mem['h0A6B]=8'h46;
    mem['h0A6C]=8'h89; mem['h0A6D]=8'h03; mem['h0A6E]=8'h26; mem['h0A6F]=8'h38;
    mem['h0A70]=8'h46; mem['h0A71]=8'hA5; mem['h0A72]=8'h02; mem['h0A73]=8'h46;
    mem['h0A74]=8'hA5; mem['h0A75]=8'h02; mem['h0A76]=8'h46; mem['h0A77]=8'h89;
    mem['h0A78]=8'h03; mem['h0A79]=8'h26; mem['h0A7A]=8'h3A; mem['h0A7B]=8'h46;
    mem['h0A7C]=8'hA5; mem['h0A7D]=8'h02; mem['h0A7E]=8'h46; mem['h0A7F]=8'hA5;
    mem['h0A80]=8'h02; mem['h0A81]=8'h46; mem['h0A82]=8'h89; mem['h0A83]=8'h03;
    mem['h0A84]=8'h44; mem['h0A85]=8'h21; mem['h0A86]=8'h0A; mem['h0A87]=8'h46;
    mem['h0A88]=8'h7E; mem['h0A89]=8'h01; mem['h0A8A]=8'h46; mem['h0A8B]=8'hDE;
    mem['h0A8C]=8'h01; mem['h0A8D]=8'h1E; mem['h0A8E]=8'h00; mem['h0A8F]=8'h46;
    mem['h0A90]=8'h20; mem['h0A91]=8'h03; mem['h0A92]=8'hA0; mem['h0A93]=8'h48;
    mem['h0A94]=8'hA5; mem['h0A95]=8'h0A; mem['h0A96]=8'h2E; mem['h0A97]=8'h38;
    mem['h0A98]=8'h2E; mem['h0A99]=8'h38; mem['h0A9A]=8'h36; mem['h0A9B]=8'h6E;
    mem['h0A9C]=8'h3E; mem['h0A9D]=8'h5D; mem['h0A9E]=8'h30; mem['h0A9F]=8'h3E;
    mem['h0AA0]=8'h01; mem['h0AA1]=8'h31; mem['h0AA2]=8'h44; mem['h0AA3]=8'hD8;
    mem['h0AA4]=8'h07; mem['h0AA5]=8'h26; mem['h0AA6]=8'h3E; mem['h0AA7]=8'h0E;
    mem['h0AA8]=8'h0A; mem['h0AA9]=8'h16; mem['h0AAA]=8'hAE; mem['h0AAB]=8'h44;
    mem['h0AAC]=8'hA9; mem['h0AAD]=8'h0B; mem['h0AAE]=8'h06; mem['h0AAF]=8'h3E;
    mem['h0AB0]=8'h46; mem['h0AB1]=8'h2C; mem['h0AB2]=8'h02; mem['h0AB3]=8'h1E;
    mem['h0AB4]=8'h00; mem['h0AB5]=8'h46; mem['h0AB6]=8'h20; mem['h0AB7]=8'h03;
    mem['h0AB8]=8'hA0; mem['h0AB9]=8'h68; mem['h0ABA]=8'h30; mem['h0ABB]=8'h0B;
    mem['h0ABC]=8'h46; mem['h0ABD]=8'h99; mem['h0ABE]=8'h02; mem['h0ABF]=8'h3C;
    mem['h0AC0]=8'h29; mem['h0AC1]=8'h68; mem['h0AC2]=8'h30; mem['h0AC3]=8'h0B;
    mem['h0AC4]=8'h3C; mem['h0AC5]=8'h20; mem['h0AC6]=8'h68; mem['h0AC7]=8'h30;
    mem['h0AC8]=8'h0B; mem['h0AC9]=8'h46; mem['h0ACA]=8'hB0; mem['h0ACB]=8'h01;
    mem['h0ACC]=8'h0E; mem['h0ACD]=8'h0A; mem['h0ACE]=8'h16; mem['h0ACF]=8'hD5;
    mem['h0AD0]=8'h26; mem['h0AD1]=8'h40; mem['h0AD2]=8'h44; mem['h0AD3]=8'hA9;
    mem['h0AD4]=8'h0B; mem['h0AD5]=8'h46; mem['h0AD6]=8'hEE; mem['h0AD7]=8'h01;
    mem['h0AD8]=8'hC8; mem['h0AD9]=8'h1E; mem['h0ADA]=8'h3E; mem['h0ADB]=8'h26;
    mem['h0ADC]=8'h40; mem['h0ADD]=8'hC3; mem['h0ADE]=8'h46; mem['h0ADF]=8'h42;
    mem['h0AE0]=8'h02; mem['h0AE1]=8'hC1; mem['h0AE2]=8'h3C; mem['h0AE3]=8'h2B;
    mem['h0AE4]=8'h68; mem['h0AE5]=8'h42; mem['h0AE6]=8'h0B; mem['h0AE7]=8'h3C;
    mem['h0AE8]=8'h2D; mem['h0AE9]=8'h68; mem['h0AEA]=8'h48; mem['h0AEB]=8'h0B;
    mem['h0AEC]=8'h3C; mem['h0AED]=8'h2A; mem['h0AEE]=8'h68; mem['h0AEF]=8'h4E;
    mem['h0AF0]=8'h0B; mem['h0AF1]=8'h3C; mem['h0AF2]=8'h2F; mem['h0AF3]=8'h68;
    mem['h0AF4]=8'h54; mem['h0AF5]=8'h0B; mem['h0AF6]=8'h3C; mem['h0AF7]=8'h3D;
    mem['h0AF8]=8'h68; mem['h0AF9]=8'h5A; mem['h0AFA]=8'h0B; mem['h0AFB]=8'h3C;
    mem['h0AFC]=8'h3C; mem['h0AFD]=8'h68; mem['h0AFE]=8'h71; mem['h0AFF]=8'h0B;
    mem['h0B00]=8'h3C; mem['h0B01]=8'h3E; mem['h0B02]=8'h68; mem['h0B03]=8'h7A;
    mem['h0B04]=8'h0B; mem['h0B05]=8'h3C; mem['h0B06]=8'h23; mem['h0B07]=8'h68;
    mem['h0B08]=8'h83; mem['h0B09]=8'h0B; mem['h0B0A]=8'h3C; mem['h0B0B]=8'h25;
    mem['h0B0C]=8'h68; mem['h0B0D]=8'h8C; mem['h0B0E]=8'h0B; mem['h0B0F]=8'h3C;
    mem['h0B10]=8'h5E; mem['h0B11]=8'h68; mem['h0B12]=8'h97; mem['h0B13]=8'h0B;
    mem['h0B14]=8'h3C; mem['h0B15]=8'h26; mem['h0B16]=8'h68; mem['h0B17]=8'h9D;
    mem['h0B18]=8'h0B; mem['h0B19]=8'h3C; mem['h0B1A]=8'h7C; mem['h0B1B]=8'h68;
    mem['h0B1C]=8'hA3; mem['h0B1D]=8'h0B; mem['h0B1E]=8'h2E; mem['h0B1F]=8'h38;
    mem['h0B20]=8'h36; mem['h0B21]=8'h70; mem['h0B22]=8'hF8; mem['h0B23]=8'h2E;
    mem['h0B24]=8'h38; mem['h0B25]=8'h36; mem['h0B26]=8'h6E; mem['h0B27]=8'h3E;
    mem['h0B28]=8'h57; mem['h0B29]=8'h30; mem['h0B2A]=8'h3E; mem['h0B2B]=8'h01;
    mem['h0B2C]=8'h31; mem['h0B2D]=8'h44; mem['h0B2E]=8'hD8; mem['h0B2F]=8'h07;
    mem['h0B30]=8'h06; mem['h0B31]=8'h52; mem['h0B32]=8'h46; mem['h0B33]=8'h42;
    mem['h0B34]=8'h02; mem['h0B35]=8'h46; mem['h0B36]=8'h1C; mem['h0B37]=8'h02;
    mem['h0B38]=8'h1E; mem['h0B39]=8'h52; mem['h0B3A]=8'h46; mem['h0B3B]=8'h65;
    mem['h0B3C]=8'h02; mem['h0B3D]=8'h1E; mem['h0B3E]=8'h00; mem['h0B3F]=8'h44;
    mem['h0B40]=8'h8E; mem['h0B41]=8'h01; mem['h0B42]=8'h46; mem['h0B43]=8'h6D;
    mem['h0B44]=8'h05; mem['h0B45]=8'h44; mem['h0B46]=8'hAE; mem['h0B47]=8'h0A;
    mem['h0B48]=8'h46; mem['h0B49]=8'h81; mem['h0B4A]=8'h05; mem['h0B4B]=8'h44;
    mem['h0B4C]=8'hAE; mem['h0B4D]=8'h0A; mem['h0B4E]=8'h46; mem['h0B4F]=8'hB5;
    mem['h0B50]=8'h05; mem['h0B51]=8'h44; mem['h0B52]=8'hAE; mem['h0B53]=8'h0A;
    mem['h0B54]=8'h46; mem['h0B55]=8'h72; mem['h0B56]=8'h06; mem['h0B57]=8'h44;
    mem['h0B58]=8'hAE; mem['h0B59]=8'h0A; mem['h0B5A]=8'h46; mem['h0B5B]=8'hFC;
    mem['h0B5C]=8'h06; mem['h0B5D]=8'h68; mem['h0B5E]=8'h66; mem['h0B5F]=8'h0B;
    mem['h0B60]=8'h46; mem['h0B61]=8'h09; mem['h0B62]=8'h05; mem['h0B63]=8'h44;
    mem['h0B64]=8'hAE; mem['h0B65]=8'h0A; mem['h0B66]=8'h2E; mem['h0B67]=8'h38;
    mem['h0B68]=8'hF3; mem['h0B69]=8'h3E; mem['h0B6A]=8'h01; mem['h0B6B]=8'h30;
    mem['h0B6C]=8'h3E; mem['h0B6D]=8'h00; mem['h0B6E]=8'h44; mem['h0B6F]=8'hAE;
    mem['h0B70]=8'h0A; mem['h0B71]=8'h46; mem['h0B72]=8'h0A; mem['h0B73]=8'h07;
    mem['h0B74]=8'h60; mem['h0B75]=8'h66; mem['h0B76]=8'h0B; mem['h0B77]=8'h44;
    mem['h0B78]=8'h60; mem['h0B79]=8'h0B; mem['h0B7A]=8'h46; mem['h0B7B]=8'h0A;
    mem['h0B7C]=8'h07; mem['h0B7D]=8'h60; mem['h0B7E]=8'h60; mem['h0B7F]=8'h0B;
    mem['h0B80]=8'h44; mem['h0B81]=8'h66; mem['h0B82]=8'h0B; mem['h0B83]=8'h46;
    mem['h0B84]=8'hFC; mem['h0B85]=8'h06; mem['h0B86]=8'h48; mem['h0B87]=8'h66;
    mem['h0B88]=8'h0B; mem['h0B89]=8'h44; mem['h0B8A]=8'h60; mem['h0B8B]=8'h0B;
    mem['h0B8C]=8'h46; mem['h0B8D]=8'h72; mem['h0B8E]=8'h06; mem['h0B8F]=8'h26;
    mem['h0B90]=8'h46; mem['h0B91]=8'h46; mem['h0B92]=8'h58; mem['h0B93]=8'h02;
    mem['h0B94]=8'h44; mem['h0B95]=8'hAE; mem['h0B96]=8'h0A; mem['h0B97]=8'h46;
    mem['h0B98]=8'hCF; mem['h0B99]=8'h06; mem['h0B9A]=8'h44; mem['h0B9B]=8'hAE;
    mem['h0B9C]=8'h0A; mem['h0B9D]=8'h46; mem['h0B9E]=8'hDE; mem['h0B9F]=8'h06;
    mem['h0BA0]=8'h44; mem['h0BA1]=8'hAE; mem['h0BA2]=8'h0A; mem['h0BA3]=8'h46;
    mem['h0BA4]=8'hED; mem['h0BA5]=8'h06; mem['h0BA6]=8'h44; mem['h0BA7]=8'hAE;
    mem['h0BA8]=8'h0A; mem['h0BA9]=8'h46; mem['h0BAA]=8'h7E; mem['h0BAB]=8'h01;
    mem['h0BAC]=8'h46; mem['h0BAD]=8'hDE; mem['h0BAE]=8'h01; mem['h0BAF]=8'h1E;
    mem['h0BB0]=8'h00; mem['h0BB1]=8'h46; mem['h0BB2]=8'h20; mem['h0BB3]=8'h03;
    mem['h0BB4]=8'h3C; mem['h0BB5]=8'h28; mem['h0BB6]=8'h68; mem['h0BB7]=8'h13;
    mem['h0BB8]=8'h0C; mem['h0BB9]=8'h26; mem['h0BBA]=8'h42; mem['h0BBB]=8'h3C;
    mem['h0BBC]=8'h2D; mem['h0BBD]=8'h68; mem['h0BBE]=8'h22; mem['h0BBF]=8'h0C;
    mem['h0BC0]=8'h46; mem['h0BC1]=8'hE0; mem['h0BC2]=8'h02; mem['h0BC3]=8'h60;
    mem['h0BC4]=8'h36; mem['h0BC5]=8'h0C; mem['h0BC6]=8'h46; mem['h0BC7]=8'h04;
    mem['h0BC8]=8'h03; mem['h0BC9]=8'h60; mem['h0BCA]=8'h3E; mem['h0BCB]=8'h0C;
    mem['h0BCC]=8'h3C; mem['h0BCD]=8'h40; mem['h0BCE]=8'h68; mem['h0BCF]=8'h4A;
    mem['h0BD0]=8'h0C; mem['h0BD1]=8'h3C; mem['h0BD2]=8'h25; mem['h0BD3]=8'h68;
    mem['h0BD4]=8'h75; mem['h0BD5]=8'h0C; mem['h0BD6]=8'h3C; mem['h0BD7]=8'h23;
    mem['h0BD8]=8'h68; mem['h0BD9]=8'h7D; mem['h0BDA]=8'h0C; mem['h0BDB]=8'h3C;
    mem['h0BDC]=8'h27; mem['h0BDD]=8'h68; mem['h0BDE]=8'h85; mem['h0BDF]=8'h0C;
    mem['h0BE0]=8'h3C; mem['h0BE1]=8'h26; mem['h0BE2]=8'h68; mem['h0BE3]=8'h98;
    mem['h0BE4]=8'h0C; mem['h0BE5]=8'h3C; mem['h0BE6]=8'h24; mem['h0BE7]=8'h68;
    mem['h0BE8]=8'hA0; mem['h0BE9]=8'h0C; mem['h0BEA]=8'h3C; mem['h0BEB]=8'h3F;
    mem['h0BEC]=8'h68; mem['h0BED]=8'hAE; mem['h0BEE]=8'h0C; mem['h0BEF]=8'h2E;
    mem['h0BF0]=8'h38; mem['h0BF1]=8'h36; mem['h0BF2]=8'h70; mem['h0BF3]=8'hF8;
    mem['h0BF4]=8'h2E; mem['h0BF5]=8'h38; mem['h0BF6]=8'h36; mem['h0BF7]=8'h6E;
    mem['h0BF8]=8'h3E; mem['h0BF9]=8'h64; mem['h0BFA]=8'h30; mem['h0BFB]=8'h3E;
    mem['h0BFC]=8'h01; mem['h0BFD]=8'h31; mem['h0BFE]=8'h44; mem['h0BFF]=8'hD8;
    mem['h0C00]=8'h07; mem['h0C01]=8'h1E; mem['h0C02]=8'h00; mem['h0C03]=8'h46;
    mem['h0C04]=8'h99; mem['h0C05]=8'h02; mem['h0C06]=8'h46; mem['h0C07]=8'h1C;
    mem['h0C08]=8'h02; mem['h0C09]=8'h1E; mem['h0C0A]=8'h42; mem['h0C0B]=8'h46;
    mem['h0C0C]=8'h65; mem['h0C0D]=8'h02; mem['h0C0E]=8'h1E; mem['h0C0F]=8'h00;
    mem['h0C10]=8'h44; mem['h0C11]=8'h8E; mem['h0C12]=8'h01; mem['h0C13]=8'h46;
    mem['h0C14]=8'h99; mem['h0C15]=8'h02; mem['h0C16]=8'h0E; mem['h0C17]=8'h0C;
    mem['h0C18]=8'h16; mem['h0C19]=8'h1F; mem['h0C1A]=8'h26; mem['h0C1B]=8'h42;
    mem['h0C1C]=8'h44; mem['h0C1D]=8'h87; mem['h0C1E]=8'h0A; mem['h0C1F]=8'h44;
    mem['h0C20]=8'h06; mem['h0C21]=8'h0C; mem['h0C22]=8'h46; mem['h0C23]=8'h99;
    mem['h0C24]=8'h02; mem['h0C25]=8'h0E; mem['h0C26]=8'h0C; mem['h0C27]=8'h16;
    mem['h0C28]=8'h2E; mem['h0C29]=8'h26; mem['h0C2A]=8'h42; mem['h0C2B]=8'h44;
    mem['h0C2C]=8'hA9; mem['h0C2D]=8'h0B; mem['h0C2E]=8'h1E; mem['h0C2F]=8'h42;
    mem['h0C30]=8'h46; mem['h0C31]=8'h48; mem['h0C32]=8'h05; mem['h0C33]=8'h44;
    mem['h0C34]=8'h06; mem['h0C35]=8'h0C; mem['h0C36]=8'h26; mem['h0C37]=8'h42;
    mem['h0C38]=8'h46; mem['h0C39]=8'h31; mem['h0C3A]=8'h04; mem['h0C3B]=8'h44;
    mem['h0C3C]=8'h06; mem['h0C3D]=8'h0C; mem['h0C3E]=8'h46; mem['h0C3F]=8'h23;
    mem['h0C40]=8'h05; mem['h0C41]=8'hE0; mem['h0C42]=8'h1E; mem['h0C43]=8'h42;
    mem['h0C44]=8'h46; mem['h0C45]=8'h58; mem['h0C46]=8'h02; mem['h0C47]=8'h44;
    mem['h0C48]=8'h01; mem['h0C49]=8'h0C; mem['h0C4A]=8'h46; mem['h0C4B]=8'h99;
    mem['h0C4C]=8'h02; mem['h0C4D]=8'h0E; mem['h0C4E]=8'h0C; mem['h0C4F]=8'h16;
    mem['h0C50]=8'h56; mem['h0C51]=8'h26; mem['h0C52]=8'h50; mem['h0C53]=8'h44;
    mem['h0C54]=8'hA9; mem['h0C55]=8'h0B; mem['h0C56]=8'hC4; mem['h0C57]=8'h46;
    mem['h0C58]=8'h99; mem['h0C59]=8'h05; mem['h0C5A]=8'h1E; mem['h0C5B]=8'h52;
    mem['h0C5C]=8'h2E; mem['h0C5D]=8'h38; mem['h0C5E]=8'hF3; mem['h0C5F]=8'h3E;
    mem['h0C60]=8'h00; mem['h0C61]=8'h30; mem['h0C62]=8'h3E; mem['h0C63]=8'h39;
    mem['h0C64]=8'h46; mem['h0C65]=8'h6D; mem['h0C66]=8'h05; mem['h0C67]=8'h26;
    mem['h0C68]=8'h42; mem['h0C69]=8'h46; mem['h0C6A]=8'h68; mem['h0C6B]=8'h03;
    mem['h0C6C]=8'h46; mem['h0C6D]=8'h99; mem['h0C6E]=8'h02; mem['h0C6F]=8'h46;
    mem['h0C70]=8'h99; mem['h0C71]=8'h02; mem['h0C72]=8'h44; mem['h0C73]=8'h06;
    mem['h0C74]=8'h0C; mem['h0C75]=8'h1E; mem['h0C76]=8'h46; mem['h0C77]=8'h46;
    mem['h0C78]=8'h65; mem['h0C79]=8'h02; mem['h0C7A]=8'h44; mem['h0C7B]=8'h01;
    mem['h0C7C]=8'h0C; mem['h0C7D]=8'h1E; mem['h0C7E]=8'h38; mem['h0C7F]=8'h46;
    mem['h0C80]=8'h65; mem['h0C81]=8'h02; mem['h0C82]=8'h44; mem['h0C83]=8'h01;
    mem['h0C84]=8'h0C; mem['h0C85]=8'h46; mem['h0C86]=8'h37; mem['h0C87]=8'h07;
    mem['h0C88]=8'h1E; mem['h0C89]=8'h4C; mem['h0C8A]=8'h46; mem['h0C8B]=8'h65;
    mem['h0C8C]=8'h02; mem['h0C8D]=8'h2E; mem['h0C8E]=8'h38; mem['h0C8F]=8'hF4;
    mem['h0C90]=8'h30; mem['h0C91]=8'hC7; mem['h0C92]=8'h24; mem['h0C93]=8'h7F;
    mem['h0C94]=8'hF8; mem['h0C95]=8'h44; mem['h0C96]=8'h01; mem['h0C97]=8'h0C;
    mem['h0C98]=8'h1E; mem['h0C99]=8'h3C; mem['h0C9A]=8'h46; mem['h0C9B]=8'h65;
    mem['h0C9C]=8'h02; mem['h0C9D]=8'h44; mem['h0C9E]=8'h01; mem['h0C9F]=8'h0C;
    mem['h0CA0]=8'h46; mem['h0CA1]=8'h4A; mem['h0CA2]=8'h00; mem['h0CA3]=8'h2E;
    mem['h0CA4]=8'h38; mem['h0CA5]=8'h36; mem['h0CA6]=8'h42; mem['h0CA7]=8'hF8;
    mem['h0CA8]=8'h30; mem['h0CA9]=8'h3E; mem['h0CAA]=8'h00; mem['h0CAB]=8'h44;
    mem['h0CAC]=8'h01; mem['h0CAD]=8'h0C; mem['h0CAE]=8'h1E; mem['h0CAF]=8'h00;
    mem['h0CB0]=8'hC3; mem['h0CB1]=8'h46; mem['h0CB2]=8'h2C; mem['h0CB3]=8'h02;
    mem['h0CB4]=8'h2E; mem['h0CB5]=8'h38; mem['h0CB6]=8'hF3; mem['h0CB7]=8'h3E;
    mem['h0CB8]=8'h00; mem['h0CB9]=8'h30; mem['h0CBA]=8'h3E; mem['h0CBB]=8'h3D;
    mem['h0CBC]=8'h46; mem['h0CBD]=8'hA8; mem['h0CBE]=8'h03; mem['h0CBF]=8'h26;
    mem['h0CC0]=8'h42; mem['h0CC1]=8'h0E; mem['h0CC2]=8'h0C; mem['h0CC3]=8'h16;
    mem['h0CC4]=8'hC8; mem['h0CC5]=8'h44; mem['h0CC6]=8'h87; mem['h0CC7]=8'h0A;
    mem['h0CC8]=8'h06; mem['h0CC9]=8'h00; mem['h0CCA]=8'h46; mem['h0CCB]=8'h42;
    mem['h0CCC]=8'h02; mem['h0CCD]=8'h44; mem['h0CCE]=8'h01; mem['h0CCF]=8'h0C;
    mem['h0CD0]=8'h1E; mem['h0CD1]=8'h00; mem['h0CD2]=8'h26; mem['h0CD3]=8'h52;
    mem['h0CD4]=8'h46; mem['h0CD5]=8'h31; mem['h0CD6]=8'h04; mem['h0CD7]=8'hF4;
    mem['h0CD8]=8'h46; mem['h0CD9]=8'h58; mem['h0CDA]=8'h05; mem['h0CDB]=8'h68;
    mem['h0CDC]=8'h24; mem['h0CDD]=8'h0D; mem['h0CDE]=8'h46; mem['h0CDF]=8'h99;
    mem['h0CE0]=8'h02; mem['h0CE1]=8'h1E; mem['h0CE2]=8'h3C; mem['h0CE3]=8'h46;
    mem['h0CE4]=8'h89; mem['h0CE5]=8'h03; mem['h0CE6]=8'h46; mem['h0CE7]=8'h99;
    mem['h0CE8]=8'h02; mem['h0CE9]=8'h46; mem['h0CEA]=8'h99; mem['h0CEB]=8'h02;
    mem['h0CEC]=8'hC3; mem['h0CED]=8'h46; mem['h0CEE]=8'h2C; mem['h0CEF]=8'h02;
    mem['h0CF0]=8'h46; mem['h0CF1]=8'h99; mem['h0CF2]=8'h02; mem['h0CF3]=8'h46;
    mem['h0CF4]=8'h99; mem['h0CF5]=8'h02; mem['h0CF6]=8'h1E; mem['h0CF7]=8'h00;
    mem['h0CF8]=8'h46; mem['h0CF9]=8'h20; mem['h0CFA]=8'h03; mem['h0CFB]=8'hA0;
    mem['h0CFC]=8'h68; mem['h0CFD]=8'h0D; mem['h0CFE]=8'h0D; mem['h0CFF]=8'h46;
    mem['h0D00]=8'h99; mem['h0D01]=8'h02; mem['h0D02]=8'h1E; mem['h0D03]=8'h3C;
    mem['h0D04]=8'h46; mem['h0D05]=8'h2F; mem['h0D06]=8'h03; mem['h0D07]=8'h46;
    mem['h0D08]=8'h99; mem['h0D09]=8'h02; mem['h0D0A]=8'h44; mem['h0D0B]=8'hF6;
    mem['h0D0C]=8'h0C; mem['h0D0D]=8'h1E; mem['h0D0E]=8'h3C; mem['h0D0F]=8'hA8;
    mem['h0D10]=8'h46; mem['h0D11]=8'h2F; mem['h0D12]=8'h03; mem['h0D13]=8'h46;
    mem['h0D14]=8'h99; mem['h0D15]=8'h02; mem['h0D16]=8'h1E; mem['h0D17]=8'h52;
    mem['h0D18]=8'hC3; mem['h0D19]=8'h46; mem['h0D1A]=8'h42; mem['h0D1B]=8'h02;
    mem['h0D1C]=8'h26; mem['h0D1D]=8'h3C; mem['h0D1E]=8'h46; mem['h0D1F]=8'h89;
    mem['h0D20]=8'h03; mem['h0D21]=8'h44; mem['h0D22]=8'h79; mem['h0D23]=8'h08;
    mem['h0D24]=8'h2E; mem['h0D25]=8'h38; mem['h0D26]=8'h36; mem['h0D27]=8'h00;
    mem['h0D28]=8'h3E; mem['h0D29]=8'h00; mem['h0D2A]=8'h30; mem['h0D2B]=8'h3E;
    mem['h0D2C]=8'h10; mem['h0D2D]=8'h31; mem['h0D2E]=8'hDE; mem['h0D2F]=8'h26;
    mem['h0D30]=8'h3C; mem['h0D31]=8'h46; mem['h0D32]=8'hFC; mem['h0D33]=8'h06;
    mem['h0D34]=8'h40; mem['h0D35]=8'hD8; mem['h0D36]=8'h07; mem['h0D37]=8'h26;
    mem['h0D38]=8'h36; mem['h0D39]=8'h46; mem['h0D3A]=8'h68; mem['h0D3B]=8'h03;
    mem['h0D3C]=8'h46; mem['h0D3D]=8'h99; mem['h0D3E]=8'h02; mem['h0D3F]=8'h46;
    mem['h0D40]=8'h99; mem['h0D41]=8'h02; mem['h0D42]=8'h46; mem['h0D43]=8'h5C;
    mem['h0D44]=8'h0D; mem['h0D45]=8'h06; mem['h0D46]=8'h20; mem['h0D47]=8'h46;
    mem['h0D48]=8'h40; mem['h0D49]=8'h00; mem['h0D4A]=8'h46; mem['h0D4B]=8'h99;
    mem['h0D4C]=8'h02; mem['h0D4D]=8'h46; mem['h0D4E]=8'h99; mem['h0D4F]=8'h02;
    mem['h0D50]=8'h46; mem['h0D51]=8'h94; mem['h0D52]=8'h0E; mem['h0D53]=8'h46;
    mem['h0D54]=8'h60; mem['h0D55]=8'h00; mem['h0D56]=8'h46; mem['h0D57]=8'h99;
    mem['h0D58]=8'h02; mem['h0D59]=8'h44; mem['h0D5A]=8'h2F; mem['h0D5B]=8'h0D;
    mem['h0D5C]=8'h46; mem['h0D5D]=8'hCE; mem['h0D5E]=8'h01; mem['h0D5F]=8'h46;
    mem['h0D60]=8'hDE; mem['h0D61]=8'h01; mem['h0D62]=8'hDC; mem['h0D63]=8'h44;
    mem['h0D64]=8'h6C; mem['h0D65]=8'h0D; mem['h0D66]=8'h46; mem['h0D67]=8'hCE;
    mem['h0D68]=8'h01; mem['h0D69]=8'h46; mem['h0D6A]=8'hDE; mem['h0D6B]=8'h01;
    mem['h0D6C]=8'h0E; mem['h0D6D]=8'h5E; mem['h0D6E]=8'h46; mem['h0D6F]=8'h72;
    mem['h0D70]=8'h02; mem['h0D71]=8'hD9; mem['h0D72]=8'h06; mem['h0D73]=8'h46;
    mem['h0D74]=8'h46; mem['h0D75]=8'h2C; mem['h0D76]=8'h02; mem['h0D77]=8'h2E;
    mem['h0D78]=8'h38; mem['h0D79]=8'h36; mem['h0D7A]=8'h73; mem['h0D7B]=8'h3E;
    mem['h0D7C]=8'h01; mem['h0D7D]=8'h46; mem['h0D7E]=8'h41; mem['h0D7F]=8'h05;
    mem['h0D80]=8'h40; mem['h0D81]=8'h8B; mem['h0D82]=8'h0D; mem['h0D83]=8'h46;
    mem['h0D84]=8'h48; mem['h0D85]=8'h05; mem['h0D86]=8'h06; mem['h0D87]=8'h2D;
    mem['h0D88]=8'h46; mem['h0D89]=8'h40; mem['h0D8A]=8'h00; mem['h0D8B]=8'h26;
    mem['h0D8C]=8'h74; mem['h0D8D]=8'h46; mem['h0D8E]=8'hEB; mem['h0D8F]=8'h05;
    mem['h0D90]=8'h46; mem['h0D91]=8'hCF; mem['h0D92]=8'h0D; mem['h0D93]=8'h26;
    mem['h0D94]=8'h46; mem['h0D95]=8'h46; mem['h0D96]=8'h58; mem['h0D97]=8'h02;
    mem['h0D98]=8'h26; mem['h0D99]=8'h76; mem['h0D9A]=8'h46; mem['h0D9B]=8'hEB;
    mem['h0D9C]=8'h05; mem['h0D9D]=8'h46; mem['h0D9E]=8'hCF; mem['h0D9F]=8'h0D;
    mem['h0DA0]=8'h26; mem['h0DA1]=8'h46; mem['h0DA2]=8'h46; mem['h0DA3]=8'h58;
    mem['h0DA4]=8'h02; mem['h0DA5]=8'h26; mem['h0DA6]=8'h78; mem['h0DA7]=8'h46;
    mem['h0DA8]=8'hEB; mem['h0DA9]=8'h05; mem['h0DAA]=8'h46; mem['h0DAB]=8'hCF;
    mem['h0DAC]=8'h0D; mem['h0DAD]=8'h26; mem['h0DAE]=8'h46; mem['h0DAF]=8'h46;
    mem['h0DB0]=8'h58; mem['h0DB1]=8'h02; mem['h0DB2]=8'h26; mem['h0DB3]=8'h7A;
    mem['h0DB4]=8'h46; mem['h0DB5]=8'hEB; mem['h0DB6]=8'h05; mem['h0DB7]=8'h46;
    mem['h0DB8]=8'hCF; mem['h0DB9]=8'h0D; mem['h0DBA]=8'h26; mem['h0DBB]=8'h46;
    mem['h0DBC]=8'h46; mem['h0DBD]=8'h58; mem['h0DBE]=8'h02; mem['h0DBF]=8'hF3;
    mem['h0DC0]=8'hC7; mem['h0DC1]=8'h46; mem['h0DC2]=8'hE3; mem['h0DC3]=8'h0D;
    mem['h0DC4]=8'h06; mem['h0DC5]=8'h46; mem['h0DC6]=8'h46; mem['h0DC7]=8'h42;
    mem['h0DC8]=8'h02; mem['h0DC9]=8'h46; mem['h0DCA]=8'h1C; mem['h0DCB]=8'h02;
    mem['h0DCC]=8'h44; mem['h0DCD]=8'h0C; mem['h0DCE]=8'h02; mem['h0DCF]=8'h2E;
    mem['h0DD0]=8'h38; mem['h0DD1]=8'hF3; mem['h0DD2]=8'hC7; mem['h0DD3]=8'h24;
    mem['h0DD4]=8'h0F; mem['h0DD5]=8'h48; mem['h0DD6]=8'hDD; mem['h0DD7]=8'h0D;
    mem['h0DD8]=8'h36; mem['h0DD9]=8'h73; mem['h0DDA]=8'hC7; mem['h0DDB]=8'hA0;
    mem['h0DDC]=8'h0B; mem['h0DDD]=8'h2E; mem['h0DDE]=8'h38; mem['h0DDF]=8'h36;
    mem['h0DE0]=8'h73; mem['h0DE1]=8'h3E; mem['h0DE2]=8'h00; mem['h0DE3]=8'h04;
    mem['h0DE4]=8'h30; mem['h0DE5]=8'h44; mem['h0DE6]=8'h40; mem['h0DE7]=8'h00;
    mem['h0DE8]=8'h2E; mem['h0DE9]=8'h38; mem['h0DEA]=8'hF3; mem['h0DEB]=8'h30;
    mem['h0DEC]=8'hC7; mem['h0DED]=8'h46; mem['h0DEE]=8'hB8; mem['h0DEF]=8'h02;
    mem['h0DF0]=8'h2E; mem['h0DF1]=8'h38; mem['h0DF2]=8'hF3; mem['h0DF3]=8'hC7;
    mem['h0DF4]=8'h44; mem['h0DF5]=8'hB8; mem['h0DF6]=8'h02; mem['h0DF7]=8'h2E;
    mem['h0DF8]=8'h38; mem['h0DF9]=8'hF4; mem['h0DFA]=8'h30; mem['h0DFB]=8'hC7;
    mem['h0DFC]=8'h46; mem['h0DFD]=8'hB8; mem['h0DFE]=8'h02; mem['h0DFF]=8'h2E;
    mem['h0E00]=8'h38; mem['h0E01]=8'hF4; mem['h0E02]=8'hC7; mem['h0E03]=8'h44;
    mem['h0E04]=8'hB8; mem['h0E05]=8'h02; mem['h0E06]=8'h46; mem['h0E07]=8'h20;
    mem['h0E08]=8'h03; mem['h0E09]=8'h3C; mem['h0E0A]=8'h3D; mem['h0E0B]=8'h48;
    mem['h0E0C]=8'hCB; mem['h0E0D]=8'h09; mem['h0E0E]=8'h46; mem['h0E0F]=8'h99;
    mem['h0E10]=8'h02; mem['h0E11]=8'h46; mem['h0E12]=8'h20; mem['h0E13]=8'h03;
    mem['h0E14]=8'hA0; mem['h0E15]=8'h68; mem['h0E16]=8'h48; mem['h0E17]=8'h0E;
    mem['h0E18]=8'h3C; mem['h0E19]=8'h22; mem['h0E1A]=8'h68; mem['h0E1B]=8'h2C;
    mem['h0E1C]=8'h0E; mem['h0E1D]=8'h26; mem['h0E1E]=8'h44; mem['h0E1F]=8'h0E;
    mem['h0E20]=8'h0E; mem['h0E21]=8'h16; mem['h0E22]=8'h26; mem['h0E23]=8'h44;
    mem['h0E24]=8'h87; mem['h0E25]=8'h0A; mem['h0E26]=8'h46; mem['h0E27]=8'h5C;
    mem['h0E28]=8'h0D; mem['h0E29]=8'h44; mem['h0E2A]=8'h4A; mem['h0E2B]=8'h09;
    mem['h0E2C]=8'h46; mem['h0E2D]=8'h99; mem['h0E2E]=8'h02; mem['h0E2F]=8'h06;
    mem['h0E30]=8'h22; mem['h0E31]=8'h46; mem['h0E32]=8'h96; mem['h0E33]=8'h0E;
    mem['h0E34]=8'h46; mem['h0E35]=8'h20; mem['h0E36]=8'h03; mem['h0E37]=8'h3C;
    mem['h0E38]=8'h3B; mem['h0E39]=8'h68; mem['h0E3A]=8'h42; mem['h0E3B]=8'h0E;
    mem['h0E3C]=8'h46; mem['h0E3D]=8'h60; mem['h0E3E]=8'h00; mem['h0E3F]=8'h44;
    mem['h0E40]=8'h4A; mem['h0E41]=8'h09; mem['h0E42]=8'h46; mem['h0E43]=8'h99;
    mem['h0E44]=8'h02; mem['h0E45]=8'h44; mem['h0E46]=8'h4A; mem['h0E47]=8'h09;
    mem['h0E48]=8'h2E; mem['h0E49]=8'h38; mem['h0E4A]=8'h36; mem['h0E4B]=8'h6E;
    mem['h0E4C]=8'h3E; mem['h0E4D]=8'h51; mem['h0E4E]=8'h30; mem['h0E4F]=8'h3E;
    mem['h0E50]=8'h01; mem['h0E51]=8'h31; mem['h0E52]=8'h44; mem['h0E53]=8'hD8;
    mem['h0E54]=8'h07; mem['h0E55]=8'h46; mem['h0E56]=8'h99; mem['h0E57]=8'h02;
    mem['h0E58]=8'h46; mem['h0E59]=8'h20; mem['h0E5A]=8'h03; mem['h0E5B]=8'h3C;
    mem['h0E5C]=8'h3D; mem['h0E5D]=8'h48; mem['h0E5E]=8'hCB; mem['h0E5F]=8'h09;
    mem['h0E60]=8'h46; mem['h0E61]=8'h99; mem['h0E62]=8'h02; mem['h0E63]=8'h26;
    mem['h0E64]=8'h44; mem['h0E65]=8'h0E; mem['h0E66]=8'h0E; mem['h0E67]=8'h16;
    mem['h0E68]=8'h6C; mem['h0E69]=8'h44; mem['h0E6A]=8'h87; mem['h0E6B]=8'h0A;
    mem['h0E6C]=8'h2E; mem['h0E6D]=8'h38; mem['h0E6E]=8'h36; mem['h0E6F]=8'h44;
    mem['h0E70]=8'hC7; mem['h0E71]=8'h46; mem['h0E72]=8'hB8; mem['h0E73]=8'h02;
    mem['h0E74]=8'h44; mem['h0E75]=8'h4A; mem['h0E76]=8'h09; mem['h0E77]=8'h46;
    mem['h0E78]=8'h99; mem['h0E79]=8'h02; mem['h0E7A]=8'h46; mem['h0E7B]=8'h20;
    mem['h0E7C]=8'h03; mem['h0E7D]=8'h3C; mem['h0E7E]=8'h3D; mem['h0E7F]=8'h48;
    mem['h0E80]=8'hCB; mem['h0E81]=8'h09; mem['h0E82]=8'h46; mem['h0E83]=8'h99;
    mem['h0E84]=8'h02; mem['h0E85]=8'h26; mem['h0E86]=8'h44; mem['h0E87]=8'h0E;
    mem['h0E88]=8'h0E; mem['h0E89]=8'h16; mem['h0E8A]=8'h8E; mem['h0E8B]=8'h44;
    mem['h0E8C]=8'h87; mem['h0E8D]=8'h0A; mem['h0E8E]=8'h46; mem['h0E8F]=8'hF7;
    mem['h0E90]=8'h0D; mem['h0E91]=8'h44; mem['h0E92]=8'h4A; mem['h0E93]=8'h09;
    mem['h0E94]=8'h06; mem['h0E95]=8'h00; mem['h0E96]=8'h46; mem['h0E97]=8'hCE;
    mem['h0E98]=8'h01; mem['h0E99]=8'h46; mem['h0E9A]=8'hDE; mem['h0E9B]=8'h01;
    mem['h0E9C]=8'hE0; mem['h0E9D]=8'h46; mem['h0E9E]=8'h3A; mem['h0E9F]=8'h05;
    mem['h0EA0]=8'hE9; mem['h0EA1]=8'hF2; mem['h0EA2]=8'h16; mem['h0EA3]=8'h00;
    mem['h0EA4]=8'hC7; mem['h0EA5]=8'hA0; mem['h0EA6]=8'h68; mem['h0EA7]=8'hBC;
    mem['h0EA8]=8'h0E; mem['h0EA9]=8'hBC; mem['h0EAA]=8'h68; mem['h0EAB]=8'hBC;
    mem['h0EAC]=8'h0E; mem['h0EAD]=8'h10; mem['h0EAE]=8'h68; mem['h0EAF]=8'hC6;
    mem['h0EB0]=8'h0E; mem['h0EB1]=8'h46; mem['h0EB2]=8'h40; mem['h0EB3]=8'h00;
    mem['h0EB4]=8'h30; mem['h0EB5]=8'h48; mem['h0EB6]=8'hA4; mem['h0EB7]=8'h0E;
    mem['h0EB8]=8'h28; mem['h0EB9]=8'h44; mem['h0EBA]=8'hA4; mem['h0EBB]=8'h0E;
    mem['h0EBC]=8'hC4; mem['h0EBD]=8'hA0; mem['h0EBE]=8'h68; mem['h0EBF]=8'hC6;
    mem['h0EC0]=8'h0E; mem['h0EC1]=8'h30; mem['h0EC2]=8'h48; mem['h0EC3]=8'hC6;
    mem['h0EC4]=8'h0E; mem['h0EC5]=8'h28; mem['h0EC6]=8'hCD; mem['h0EC7]=8'hD6;
    mem['h0EC8]=8'h46; mem['h0EC9]=8'h1C; mem['h0ECA]=8'h02; mem['h0ECB]=8'h46;
    mem['h0ECC]=8'h33; mem['h0ECD]=8'h05; mem['h0ECE]=8'h44; mem['h0ECF]=8'h0C;
    mem['h0ED0]=8'h02; mem['h0ED1]=8'h00; mem['h0ED2]=8'h00; mem['h0ED3]=8'h00;
end
