// rom.v
// to be included from the top module at the comple

initial
begin
    mem['hE000]=8'h8D; mem['hE001]=8'h03; mem['hE002]=8'h27; mem['hE003]=8'hFC;
    mem['hE004]=8'h39; mem['hE005]=8'hB6; mem['hE006]=8'h80; mem['hE007]=8'h18;
    mem['hE008]=8'h85; mem['hE009]=8'h01; mem['hE00A]=8'h27; mem['hE00B]=8'h06;
    mem['hE00C]=8'hB6; mem['hE00D]=8'h80; mem['hE00E]=8'h19; mem['hE00F]=8'h84;
    mem['hE010]=8'h7F; mem['hE011]=8'h39; mem['hE012]=8'h4F; mem['hE013]=8'h39;
    mem['hE014]=8'h8D; mem['hE015]=8'h24; mem['hE016]=8'h34; mem['hE017]=8'h02;
    mem['hE018]=8'h81; mem['hE019]=8'h0D; mem['hE01A]=8'h27; mem['hE01B]=8'h0B;
    mem['hE01C]=8'hB7; mem['hE01D]=8'h80; mem['hE01E]=8'h19; mem['hE01F]=8'h0C;
    mem['hE020]=8'h79; mem['hE021]=8'h96; mem['hE022]=8'h79; mem['hE023]=8'h91;
    mem['hE024]=8'h78; mem['hE025]=8'h25; mem['hE026]=8'h10; mem['hE027]=8'h0F;
    mem['hE028]=8'h79; mem['hE029]=8'h8D; mem['hE02A]=8'h0F; mem['hE02B]=8'h86;
    mem['hE02C]=8'h0D; mem['hE02D]=8'hB7; mem['hE02E]=8'h80; mem['hE02F]=8'h19;
    mem['hE030]=8'h8D; mem['hE031]=8'h08; mem['hE032]=8'h86; mem['hE033]=8'h0A;
    mem['hE034]=8'hB7; mem['hE035]=8'h80; mem['hE036]=8'h19; mem['hE037]=8'h35;
    mem['hE038]=8'h02; mem['hE039]=8'h39; mem['hE03A]=8'h34; mem['hE03B]=8'h02;
    mem['hE03C]=8'hB6; mem['hE03D]=8'h80; mem['hE03E]=8'h18; mem['hE03F]=8'h85;
    mem['hE040]=8'h02; mem['hE041]=8'h27; mem['hE042]=8'hF9; mem['hE043]=8'h35;
    mem['hE044]=8'h02; mem['hE045]=8'h39; mem['hE046]=8'h10; mem['hE047]=8'hCE;
    mem['hE048]=8'h01; mem['hE049]=8'hEE; mem['hE04A]=8'h96; mem['hE04B]=8'h6E;
    mem['hE04C]=8'h81; mem['hE04D]=8'h55; mem['hE04E]=8'h26; mem['hE04F]=8'h0A;
    mem['hE050]=8'h9E; mem['hE051]=8'h6F; mem['hE052]=8'hA6; mem['hE053]=8'h84;
    mem['hE054]=8'h81; mem['hE055]=8'h12; mem['hE056]=8'h26; mem['hE057]=8'h02;
    mem['hE058]=8'h6E; mem['hE059]=8'h84; mem['hE05A]=8'h8E; mem['hE05B]=8'h02;
    mem['hE05C]=8'h18; mem['hE05D]=8'h6F; mem['hE05E]=8'h83; mem['hE05F]=8'h30;
    mem['hE060]=8'h01; mem['hE061]=8'h26; mem['hE062]=8'hFA; mem['hE063]=8'h8E;
    mem['hE064]=8'h02; mem['hE065]=8'h17; mem['hE066]=8'h6F; mem['hE067]=8'h80;
    mem['hE068]=8'h9F; mem['hE069]=8'h19; mem['hE06A]=8'hA6; mem['hE06B]=8'h02;
    mem['hE06C]=8'h43; mem['hE06D]=8'hA7; mem['hE06E]=8'h02; mem['hE06F]=8'hA1;
    mem['hE070]=8'h02; mem['hE071]=8'h26; mem['hE072]=8'h06; mem['hE073]=8'h30;
    mem['hE074]=8'h01; mem['hE075]=8'h63; mem['hE076]=8'h01; mem['hE077]=8'h20;
    mem['hE078]=8'hF1; mem['hE079]=8'h9F; mem['hE07A]=8'h71; mem['hE07B]=8'h9F;
    mem['hE07C]=8'h27; mem['hE07D]=8'h9F; mem['hE07E]=8'h23; mem['hE07F]=8'h30;
    mem['hE080]=8'h89; mem['hE081]=8'hFF; mem['hE082]=8'h38; mem['hE083]=8'h9F;
    mem['hE084]=8'h21; mem['hE085]=8'h1F; mem['hE086]=8'h14; mem['hE087]=8'h8E;
    mem['hE088]=8'hE0; mem['hE089]=8'hCE; mem['hE08A]=8'hCE; mem['hE08B]=8'h00;
    mem['hE08C]=8'h76; mem['hE08D]=8'hC6; mem['hE08E]=8'h12; mem['hE08F]=8'hBD;
    mem['hE090]=8'hE1; mem['hE091]=8'hAE; mem['hE092]=8'hCE; mem['hE093]=8'h00;
    mem['hE094]=8'hA7; mem['hE095]=8'hC6; mem['hE096]=8'h04; mem['hE097]=8'hBD;
    mem['hE098]=8'hE1; mem['hE099]=8'hAE; mem['hE09A]=8'h86; mem['hE09B]=8'h39;
    mem['hE09C]=8'h97; mem['hE09D]=8'hF0; mem['hE09E]=8'hBD; mem['hE09F]=8'hE4;
    mem['hE0A0]=8'hBA; mem['hE0A1]=8'h8E; mem['hE0A2]=8'h00; mem['hE0A3]=8'hB5;
    mem['hE0A4]=8'h9F; mem['hE0A5]=8'h8D; mem['hE0A6]=8'hCE; mem['hE0A7]=8'hEB;
    mem['hE0A8]=8'hCE; mem['hE0A9]=8'hC6; mem['hE0AA]=8'h0A; mem['hE0AB]=8'hEF;
    mem['hE0AC]=8'h81; mem['hE0AD]=8'h5A; mem['hE0AE]=8'h26; mem['hE0AF]=8'hFB;
    mem['hE0B0]=8'h86; mem['hE0B1]=8'h15; mem['hE0B2]=8'hB7; mem['hE0B3]=8'h80;
    mem['hE0B4]=8'h18; mem['hE0B5]=8'h8E; mem['hE0B6]=8'hE1; mem['hE0B7]=8'h03;
    mem['hE0B8]=8'hBD; mem['hE0B9]=8'hF0; mem['hE0BA]=8'hE2; mem['hE0BB]=8'h8E;
    mem['hE0BC]=8'hE0; mem['hE0BD]=8'hC6; mem['hE0BE]=8'h9F; mem['hE0BF]=8'h6F;
    mem['hE0C0]=8'h86; mem['hE0C1]=8'h55; mem['hE0C2]=8'h97; mem['hE0C3]=8'h6E;
    mem['hE0C4]=8'h20; mem['hE0C5]=8'h04; mem['hE0C6]=8'h12; mem['hE0C7]=8'hBD;
    mem['hE0C8]=8'hE4; mem['hE0C9]=8'hD4; mem['hE0CA]=8'h7E; mem['hE0CB]=8'hE4;
    mem['hE0CC]=8'h22; mem['hE0CD]=8'h3B; mem['hE0CE]=8'h10; mem['hE0CF]=8'h40;
    mem['hE0D0]=8'hFF; mem['hE0D1]=8'h00; mem['hE0D2]=8'hEB; mem['hE0D3]=8'hCE;
    mem['hE0D4]=8'h0C; mem['hE0D5]=8'h84; mem['hE0D6]=8'h26; mem['hE0D7]=8'h02;
    mem['hE0D8]=8'h0C; mem['hE0D9]=8'h83; mem['hE0DA]=8'hB6; mem['hE0DB]=8'h00;
    mem['hE0DC]=8'h00; mem['hE0DD]=8'h7E; mem['hE0DE]=8'hE1; mem['hE0DF]=8'hBF;
    mem['hE0E0]=8'h7E; mem['hE0E1]=8'hE1; mem['hE0E2]=8'hBE; mem['hE0E3]=8'h7E;
    mem['hE0E4]=8'hE0; mem['hE0E5]=8'hCD; mem['hE0E6]=8'h7E; mem['hE0E7]=8'hEB;
    mem['hE0E8]=8'hCE; mem['hE0E9]=8'h80; mem['hE0EA]=8'h4F; mem['hE0EB]=8'hC7;
    mem['hE0EC]=8'h52; mem['hE0ED]=8'h59; mem['hE0EE]=8'h32; mem['hE0EF]=8'hE2;
    mem['hE0F0]=8'h1D; mem['hE0F1]=8'hE3; mem['hE0F2]=8'h2A; mem['hE0F3]=8'h1D;
    mem['hE0F4]=8'hE2; mem['hE0F5]=8'hBD; mem['hE0F6]=8'hE1; mem['hE0F7]=8'hCE;
    mem['hE0F8]=8'h00; mem['hE0F9]=8'h00; mem['hE0FA]=8'h00; mem['hE0FB]=8'h00;
    mem['hE0FC]=8'h00; mem['hE0FD]=8'h00; mem['hE0FE]=8'h00; mem['hE0FF]=8'h00;
    mem['hE100]=8'h00; mem['hE101]=8'h00; mem['hE102]=8'h00; mem['hE103]=8'h00;
    mem['hE104]=8'h36; mem['hE105]=8'h38; mem['hE106]=8'h30; mem['hE107]=8'h39;
    mem['hE108]=8'h20; mem['hE109]=8'h45; mem['hE10A]=8'h58; mem['hE10B]=8'h54;
    mem['hE10C]=8'h45; mem['hE10D]=8'h4E; mem['hE10E]=8'h44; mem['hE10F]=8'h45;
    mem['hE110]=8'h44; mem['hE111]=8'h20; mem['hE112]=8'h42; mem['hE113]=8'h41;
    mem['hE114]=8'h53; mem['hE115]=8'h49; mem['hE116]=8'h43; mem['hE117]=8'h0D;
    mem['hE118]=8'h28; mem['hE119]=8'h43; mem['hE11A]=8'h29; mem['hE11B]=8'h20;
    mem['hE11C]=8'h31; mem['hE11D]=8'h39; mem['hE11E]=8'h38; mem['hE11F]=8'h32;
    mem['hE120]=8'h20; mem['hE121]=8'h42; mem['hE122]=8'h59; mem['hE123]=8'h20;
    mem['hE124]=8'h4D; mem['hE125]=8'h49; mem['hE126]=8'h43; mem['hE127]=8'h52;
    mem['hE128]=8'h4F; mem['hE129]=8'h53; mem['hE12A]=8'h4F; mem['hE12B]=8'h46;
    mem['hE12C]=8'h54; mem['hE12D]=8'h0D; mem['hE12E]=8'h0D; mem['hE12F]=8'h00;
    mem['hE130]=8'h34; mem['hE131]=8'h16; mem['hE132]=8'h9E; mem['hE133]=8'h76;
    mem['hE134]=8'hDC; mem['hE135]=8'h78; mem['hE136]=8'h9F; mem['hE137]=8'h6A;
    mem['hE138]=8'hD7; mem['hE139]=8'h6C; mem['hE13A]=8'h97; mem['hE13B]=8'h6D;
    mem['hE13C]=8'h35; mem['hE13D]=8'h96; mem['hE13E]=8'h0F; mem['hE13F]=8'h73;
    mem['hE140]=8'h8E; mem['hE141]=8'h00; mem['hE142]=8'hF4; mem['hE143]=8'hC6;
    mem['hE144]=8'h01; mem['hE145]=8'hBD; mem['hE146]=8'hE0; mem['hE147]=8'h00;
    mem['hE148]=8'h81; mem['hE149]=8'h08; mem['hE14A]=8'h26; mem['hE14B]=8'h07;
    mem['hE14C]=8'h5A; mem['hE14D]=8'h27; mem['hE14E]=8'hEF; mem['hE14F]=8'h30;
    mem['hE150]=8'h1F; mem['hE151]=8'h20; mem['hE152]=8'h34; mem['hE153]=8'h81;
    mem['hE154]=8'h15; mem['hE155]=8'h26; mem['hE156]=8'h0A; mem['hE157]=8'h5A;
    mem['hE158]=8'h27; mem['hE159]=8'hE4; mem['hE15A]=8'h86; mem['hE15B]=8'h08;
    mem['hE15C]=8'hBD; mem['hE15D]=8'hE0; mem['hE15E]=8'h14; mem['hE15F]=8'h20;
    mem['hE160]=8'hF6; mem['hE161]=8'h81; mem['hE162]=8'h03; mem['hE163]=8'h1A;
    mem['hE164]=8'h01; mem['hE165]=8'h27; mem['hE166]=8'h05; mem['hE167]=8'h81;
    mem['hE168]=8'h0D; mem['hE169]=8'h26; mem['hE16A]=8'h0D; mem['hE16B]=8'h4F;
    mem['hE16C]=8'h34; mem['hE16D]=8'h01; mem['hE16E]=8'hBD; mem['hE16F]=8'hF0;
    mem['hE170]=8'hA2; mem['hE171]=8'h6F; mem['hE172]=8'h84; mem['hE173]=8'h8E;
    mem['hE174]=8'h00; mem['hE175]=8'hF3; mem['hE176]=8'h35; mem['hE177]=8'h81;
    mem['hE178]=8'h81; mem['hE179]=8'h20; mem['hE17A]=8'h25; mem['hE17B]=8'hC9;
    mem['hE17C]=8'h81; mem['hE17D]=8'h7B; mem['hE17E]=8'h24; mem['hE17F]=8'hC5;
    mem['hE180]=8'hC1; mem['hE181]=8'hFA; mem['hE182]=8'h24; mem['hE183]=8'hC1;
    mem['hE184]=8'hA7; mem['hE185]=8'h80; mem['hE186]=8'h5C; mem['hE187]=8'hBD;
    mem['hE188]=8'hE0; mem['hE189]=8'h14; mem['hE18A]=8'h20; mem['hE18B]=8'hB9;
    mem['hE18C]=8'h27; mem['hE18D]=8'h05; mem['hE18E]=8'hBD; mem['hE18F]=8'hEE;
    mem['hE190]=8'hC1; mem['hE191]=8'h9F; mem['hE192]=8'h7A; mem['hE193]=8'h6E;
    mem['hE194]=8'h9F; mem['hE195]=8'h00; mem['hE196]=8'h7A; mem['hE197]=8'h7E;
    mem['hE198]=8'hE5; mem['hE199]=8'hA3; mem['hE19A]=8'h96; mem['hE19B]=8'h73;
    mem['hE19C]=8'h26; mem['hE19D]=8'h03; mem['hE19E]=8'hBD; mem['hE19F]=8'hE0;
    mem['hE1A0]=8'h05; mem['hE1A1]=8'h0F; mem['hE1A2]=8'h73; mem['hE1A3]=8'h97;
    mem['hE1A4]=8'h53; mem['hE1A5]=8'h10; mem['hE1A6]=8'h26; mem['hE1A7]=8'h0C;
    mem['hE1A8]=8'h6A; mem['hE1A9]=8'h97; mem['hE1AA]=8'h56; mem['hE1AB]=8'h7E;
    mem['hE1AC]=8'hEE; mem['hE1AD]=8'h1F; mem['hE1AE]=8'hA6; mem['hE1AF]=8'h80;
    mem['hE1B0]=8'hA7; mem['hE1B1]=8'hC0; mem['hE1B2]=8'h5A; mem['hE1B3]=8'h26;
    mem['hE1B4]=8'hF9; mem['hE1B5]=8'h39; mem['hE1B6]=8'h39; mem['hE1B7]=8'h9D;
    mem['hE1B8]=8'h82; mem['hE1B9]=8'h27; mem['hE1BA]=8'hFB; mem['hE1BB]=8'h7E;
    mem['hE1BC]=8'hEA; mem['hE1BD]=8'h00; mem['hE1BE]=8'h3B; mem['hE1BF]=8'h81;
    mem['hE1C0]=8'h3A; mem['hE1C1]=8'h24; mem['hE1C2]=8'h0A; mem['hE1C3]=8'h81;
    mem['hE1C4]=8'h20; mem['hE1C5]=8'h26; mem['hE1C6]=8'h02; mem['hE1C7]=8'h0E;
    mem['hE1C8]=8'h7C; mem['hE1C9]=8'h80; mem['hE1CA]=8'h30; mem['hE1CB]=8'h80;
    mem['hE1CC]=8'hD0; mem['hE1CD]=8'h39; mem['hE1CE]=8'hF3; mem['hE1CF]=8'hC0;
    mem['hE1D0]=8'hF4; mem['hE1D1]=8'h34; mem['hE1D2]=8'hF3; mem['hE1D3]=8'hD9;
    mem['hE1D4]=8'h00; mem['hE1D5]=8'hAD; mem['hE1D6]=8'hF6; mem['hE1D7]=8'h65;
    mem['hE1D8]=8'hF6; mem['hE1D9]=8'hBA; mem['hE1DA]=8'hEE; mem['hE1DB]=8'hD4;
    mem['hE1DC]=8'hEE; mem['hE1DD]=8'h05; mem['hE1DE]=8'hEC; mem['hE1DF]=8'h81;
    mem['hE1E0]=8'hEE; mem['hE1E1]=8'h9A; mem['hE1E2]=8'hEE; mem['hE1E3]=8'h24;
    mem['hE1E4]=8'hEE; mem['hE1E5]=8'h10; mem['hE1E6]=8'hF7; mem['hE1E7]=8'h6A;
    mem['hE1E8]=8'hF7; mem['hE1E9]=8'h32; mem['hE1EA]=8'hF7; mem['hE1EB]=8'h3B;
    mem['hE1EC]=8'hF8; mem['hE1ED]=8'hAC; mem['hE1EE]=8'hF8; mem['hE1EF]=8'hDE;
    mem['hE1F0]=8'hF8; mem['hE1F1]=8'h00; mem['hE1F2]=8'hFA; mem['hE1F3]=8'h66;
    mem['hE1F4]=8'hF8; mem['hE1F5]=8'h3A; mem['hE1F6]=8'hFF; mem['hE1F7]=8'h38;
    mem['hE1F8]=8'hEE; mem['hE1F9]=8'h2F; mem['hE1FA]=8'hEE; mem['hE1FB]=8'h4C;
    mem['hE1FC]=8'hEE; mem['hE1FD]=8'h53; mem['hE1FE]=8'hE1; mem['hE1FF]=8'h9A;
    mem['hE200]=8'hEC; mem['hE201]=8'h72; mem['hE202]=8'hFA; mem['hE203]=8'h6E;
    mem['hE204]=8'hFB; mem['hE205]=8'h2E; mem['hE206]=8'hFA; mem['hE207]=8'hFE;
    mem['hE208]=8'h79; mem['hE209]=8'hF1; mem['hE20A]=8'h0B; mem['hE20B]=8'h79;
    mem['hE20C]=8'hF1; mem['hE20D]=8'h02; mem['hE20E]=8'h7B; mem['hE20F]=8'hF2;
    mem['hE210]=8'h12; mem['hE211]=8'h7B; mem['hE212]=8'hF2; mem['hE213]=8'hD7;
    mem['hE214]=8'h7F; mem['hE215]=8'hF8; mem['hE216]=8'h43; mem['hE217]=8'h50;
    mem['hE218]=8'hEA; mem['hE219]=8'h59; mem['hE21A]=8'h46; mem['hE21B]=8'hEA;
    mem['hE21C]=8'h58; mem['hE21D]=8'h46; mem['hE21E]=8'h4F; mem['hE21F]=8'hD2;
    mem['hE220]=8'h47; mem['hE221]=8'hCF; mem['hE222]=8'h52; mem['hE223]=8'h45;
    mem['hE224]=8'hCD; mem['hE225]=8'hA7; mem['hE226]=8'h45; mem['hE227]=8'h4C;
    mem['hE228]=8'h53; mem['hE229]=8'hC5; mem['hE22A]=8'h49; mem['hE22B]=8'hC6;
    mem['hE22C]=8'h44; mem['hE22D]=8'h41; mem['hE22E]=8'h54; mem['hE22F]=8'hC1;
    mem['hE230]=8'h50; mem['hE231]=8'h52; mem['hE232]=8'h49; mem['hE233]=8'h4E;
    mem['hE234]=8'hD4; mem['hE235]=8'h4F; mem['hE236]=8'hCE; mem['hE237]=8'h49;
    mem['hE238]=8'h4E; mem['hE239]=8'h50; mem['hE23A]=8'h55; mem['hE23B]=8'hD4;
    mem['hE23C]=8'h45; mem['hE23D]=8'h4E; mem['hE23E]=8'hC4; mem['hE23F]=8'h4E;
    mem['hE240]=8'h45; mem['hE241]=8'h58; mem['hE242]=8'hD4; mem['hE243]=8'h44;
    mem['hE244]=8'h49; mem['hE245]=8'hCD; mem['hE246]=8'h52; mem['hE247]=8'h45;
    mem['hE248]=8'h41; mem['hE249]=8'hC4; mem['hE24A]=8'h52; mem['hE24B]=8'h55;
    mem['hE24C]=8'hCE; mem['hE24D]=8'h52; mem['hE24E]=8'h45; mem['hE24F]=8'h53;
    mem['hE250]=8'h54; mem['hE251]=8'h4F; mem['hE252]=8'h52; mem['hE253]=8'hC5;
    mem['hE254]=8'h52; mem['hE255]=8'h45; mem['hE256]=8'h54; mem['hE257]=8'h55;
    mem['hE258]=8'h52; mem['hE259]=8'hCE; mem['hE25A]=8'h53; mem['hE25B]=8'h54;
    mem['hE25C]=8'h4F; mem['hE25D]=8'hD0; mem['hE25E]=8'h50; mem['hE25F]=8'h4F;
    mem['hE260]=8'h4B; mem['hE261]=8'hC5; mem['hE262]=8'h43; mem['hE263]=8'h4F;
    mem['hE264]=8'h4E; mem['hE265]=8'hD4; mem['hE266]=8'h4C; mem['hE267]=8'h49;
    mem['hE268]=8'h53; mem['hE269]=8'hD4; mem['hE26A]=8'h43; mem['hE26B]=8'h4C;
    mem['hE26C]=8'h45; mem['hE26D]=8'h41; mem['hE26E]=8'hD2; mem['hE26F]=8'h4E;
    mem['hE270]=8'h45; mem['hE271]=8'hD7; mem['hE272]=8'h45; mem['hE273]=8'h58;
    mem['hE274]=8'h45; mem['hE275]=8'hC3; mem['hE276]=8'h54; mem['hE277]=8'h52;
    mem['hE278]=8'h4F; mem['hE279]=8'hCE; mem['hE27A]=8'h54; mem['hE27B]=8'h52;
    mem['hE27C]=8'h4F; mem['hE27D]=8'h46; mem['hE27E]=8'hC6; mem['hE27F]=8'h44;
    mem['hE280]=8'h45; mem['hE281]=8'hCC; mem['hE282]=8'h44; mem['hE283]=8'h45;
    mem['hE284]=8'hC6; mem['hE285]=8'h4C; mem['hE286]=8'h49; mem['hE287]=8'h4E;
    mem['hE288]=8'hC5; mem['hE289]=8'h52; mem['hE28A]=8'h45; mem['hE28B]=8'h4E;
    mem['hE28C]=8'h55; mem['hE28D]=8'hCD; mem['hE28E]=8'h45; mem['hE28F]=8'h44;
    mem['hE290]=8'h49; mem['hE291]=8'hD4; mem['hE292]=8'h54; mem['hE293]=8'h41;
    mem['hE294]=8'h42; mem['hE295]=8'hA8; mem['hE296]=8'h54; mem['hE297]=8'hCF;
    mem['hE298]=8'h53; mem['hE299]=8'h55; mem['hE29A]=8'hC2; mem['hE29B]=8'h54;
    mem['hE29C]=8'h48; mem['hE29D]=8'h45; mem['hE29E]=8'hCE; mem['hE29F]=8'h4E;
    mem['hE2A0]=8'h4F; mem['hE2A1]=8'hD4; mem['hE2A2]=8'h53; mem['hE2A3]=8'h54;
    mem['hE2A4]=8'h45; mem['hE2A5]=8'hD0; mem['hE2A6]=8'h4F; mem['hE2A7]=8'h46;
    mem['hE2A8]=8'hC6; mem['hE2A9]=8'hAB; mem['hE2AA]=8'hAD; mem['hE2AB]=8'hAA;
    mem['hE2AC]=8'hAF; mem['hE2AD]=8'hDE; mem['hE2AE]=8'h41; mem['hE2AF]=8'h4E;
    mem['hE2B0]=8'hC4; mem['hE2B1]=8'h4F; mem['hE2B2]=8'hD2; mem['hE2B3]=8'hBE;
    mem['hE2B4]=8'hBD; mem['hE2B5]=8'hBC; mem['hE2B6]=8'h46; mem['hE2B7]=8'hCE;
    mem['hE2B8]=8'h55; mem['hE2B9]=8'h53; mem['hE2BA]=8'h49; mem['hE2BB]=8'h4E;
    mem['hE2BC]=8'hC7; mem['hE2BD]=8'h53; mem['hE2BE]=8'h47; mem['hE2BF]=8'hCE;
    mem['hE2C0]=8'h49; mem['hE2C1]=8'h4E; mem['hE2C2]=8'hD4; mem['hE2C3]=8'h41;
    mem['hE2C4]=8'h42; mem['hE2C5]=8'hD3; mem['hE2C6]=8'h55; mem['hE2C7]=8'h53;
    mem['hE2C8]=8'hD2; mem['hE2C9]=8'h52; mem['hE2CA]=8'h4E; mem['hE2CB]=8'hC4;
    mem['hE2CC]=8'h53; mem['hE2CD]=8'h49; mem['hE2CE]=8'hCE; mem['hE2CF]=8'h50;
    mem['hE2D0]=8'h45; mem['hE2D1]=8'h45; mem['hE2D2]=8'hCB; mem['hE2D3]=8'h4C;
    mem['hE2D4]=8'h45; mem['hE2D5]=8'hCE; mem['hE2D6]=8'h53; mem['hE2D7]=8'h54;
    mem['hE2D8]=8'h52; mem['hE2D9]=8'hA4; mem['hE2DA]=8'h56; mem['hE2DB]=8'h41;
    mem['hE2DC]=8'hCC; mem['hE2DD]=8'h41; mem['hE2DE]=8'h53; mem['hE2DF]=8'hC3;
    mem['hE2E0]=8'h43; mem['hE2E1]=8'h48; mem['hE2E2]=8'h52; mem['hE2E3]=8'hA4;
    mem['hE2E4]=8'h41; mem['hE2E5]=8'h54; mem['hE2E6]=8'hCE; mem['hE2E7]=8'h43;
    mem['hE2E8]=8'h4F; mem['hE2E9]=8'hD3; mem['hE2EA]=8'h54; mem['hE2EB]=8'h41;
    mem['hE2EC]=8'hCE; mem['hE2ED]=8'h45; mem['hE2EE]=8'h58; mem['hE2EF]=8'hD0;
    mem['hE2F0]=8'h46; mem['hE2F1]=8'h49; mem['hE2F2]=8'hD8; mem['hE2F3]=8'h4C;
    mem['hE2F4]=8'h4F; mem['hE2F5]=8'hC7; mem['hE2F6]=8'h50; mem['hE2F7]=8'h4F;
    mem['hE2F8]=8'hD3; mem['hE2F9]=8'h53; mem['hE2FA]=8'h51; mem['hE2FB]=8'hD2;
    mem['hE2FC]=8'h48; mem['hE2FD]=8'h45; mem['hE2FE]=8'h58; mem['hE2FF]=8'hA4;
    mem['hE300]=8'h4C; mem['hE301]=8'h45; mem['hE302]=8'h46; mem['hE303]=8'h54;
    mem['hE304]=8'hA4; mem['hE305]=8'h52; mem['hE306]=8'h49; mem['hE307]=8'h47;
    mem['hE308]=8'h48; mem['hE309]=8'h54; mem['hE30A]=8'hA4; mem['hE30B]=8'h4D;
    mem['hE30C]=8'h49; mem['hE30D]=8'h44; mem['hE30E]=8'hA4; mem['hE30F]=8'h49;
    mem['hE310]=8'h4E; mem['hE311]=8'h4B; mem['hE312]=8'h45; mem['hE313]=8'h59;
    mem['hE314]=8'hA4; mem['hE315]=8'h4D; mem['hE316]=8'h45; mem['hE317]=8'hCD;
    mem['hE318]=8'h56; mem['hE319]=8'h41; mem['hE31A]=8'h52; mem['hE31B]=8'h50;
    mem['hE31C]=8'h54; mem['hE31D]=8'hD2; mem['hE31E]=8'h49; mem['hE31F]=8'h4E;
    mem['hE320]=8'h53; mem['hE321]=8'h54; mem['hE322]=8'hD2; mem['hE323]=8'h53;
    mem['hE324]=8'h54; mem['hE325]=8'h52; mem['hE326]=8'h49; mem['hE327]=8'h4E;
    mem['hE328]=8'h47; mem['hE329]=8'hA4; mem['hE32A]=8'hE4; mem['hE32B]=8'hE8;
    mem['hE32C]=8'hE6; mem['hE32D]=8'h33; mem['hE32E]=8'hE6; mem['hE32F]=8'h90;
    mem['hE330]=8'hE6; mem['hE331]=8'h90; mem['hE332]=8'hE6; mem['hE333]=8'h90;
    mem['hE334]=8'hE6; mem['hE335]=8'hC1; mem['hE336]=8'hE6; mem['hE337]=8'h8D;
    mem['hE338]=8'hF0; mem['hE339]=8'h6A; mem['hE33A]=8'hE6; mem['hE33B]=8'hEF;
    mem['hE33C]=8'hE7; mem['hE33D]=8'h9C; mem['hE33E]=8'hE5; mem['hE33F]=8'hBA;
    mem['hE340]=8'hE8; mem['hE341]=8'h81; mem['hE342]=8'hEA; mem['hE343]=8'hD2;
    mem['hE344]=8'hE7; mem['hE345]=8'hD6; mem['hE346]=8'hE6; mem['hE347]=8'h28;
    mem['hE348]=8'hE5; mem['hE349]=8'h9C; mem['hE34A]=8'hE6; mem['hE34B]=8'h6D;
    mem['hE34C]=8'hE5; mem['hE34D]=8'hBE; mem['hE34E]=8'hEE; mem['hE34F]=8'hDB;
    mem['hE350]=8'hE5; mem['hE351]=8'hE3; mem['hE352]=8'hEE; mem['hE353]=8'hE2;
    mem['hE354]=8'hE5; mem['hE355]=8'hF4; mem['hE356]=8'hE4; mem['hE357]=8'hB8;
    mem['hE358]=8'hE1; mem['hE359]=8'h8C; mem['hE35A]=8'hFA; mem['hE35B]=8'h61;
    mem['hE35C]=8'hFA; mem['hE35D]=8'h62; mem['hE35E]=8'hFC; mem['hE35F]=8'hDD;
    mem['hE360]=8'hFC; mem['hE361]=8'h21; mem['hE362]=8'hFF; mem['hE363]=8'h7C;
    mem['hE364]=8'hFD; mem['hE365]=8'h67; mem['hE366]=8'hF8; mem['hE367]=8'hED;
    mem['hE368]=8'h4E; mem['hE369]=8'h46; mem['hE36A]=8'h53; mem['hE36B]=8'h4E;
    mem['hE36C]=8'h52; mem['hE36D]=8'h47; mem['hE36E]=8'h4F; mem['hE36F]=8'h44;
    mem['hE370]=8'h46; mem['hE371]=8'h43; mem['hE372]=8'h4F; mem['hE373]=8'h56;
    mem['hE374]=8'h4F; mem['hE375]=8'h4D; mem['hE376]=8'h55; mem['hE377]=8'h4C;
    mem['hE378]=8'h42; mem['hE379]=8'h53; mem['hE37A]=8'h44; mem['hE37B]=8'h44;
    mem['hE37C]=8'h2F; mem['hE37D]=8'h30; mem['hE37E]=8'h49; mem['hE37F]=8'h44;
    mem['hE380]=8'h54; mem['hE381]=8'h4D; mem['hE382]=8'h4F; mem['hE383]=8'h53;
    mem['hE384]=8'h4C; mem['hE385]=8'h53; mem['hE386]=8'h53; mem['hE387]=8'h54;
    mem['hE388]=8'h43; mem['hE389]=8'h4E; mem['hE38A]=8'h46; mem['hE38B]=8'h44;
    mem['hE38C]=8'h41; mem['hE38D]=8'h4F; mem['hE38E]=8'h44; mem['hE38F]=8'h4E;
    mem['hE390]=8'h49; mem['hE391]=8'h4F; mem['hE392]=8'h46; mem['hE393]=8'h4D;
    mem['hE394]=8'h4E; mem['hE395]=8'h4F; mem['hE396]=8'h49; mem['hE397]=8'h45;
    mem['hE398]=8'h44; mem['hE399]=8'h53; mem['hE39A]=8'h55; mem['hE39B]=8'h46;
    mem['hE39C]=8'h4E; mem['hE39D]=8'h45; mem['hE39E]=8'h20; mem['hE39F]=8'h45;
    mem['hE3A0]=8'h52; mem['hE3A1]=8'h52; mem['hE3A2]=8'h4F; mem['hE3A3]=8'h52;
    mem['hE3A4]=8'h00; mem['hE3A5]=8'h20; mem['hE3A6]=8'h49; mem['hE3A7]=8'h4E;
    mem['hE3A8]=8'h20; mem['hE3A9]=8'h00; mem['hE3AA]=8'h0D; mem['hE3AB]=8'h4F;
    mem['hE3AC]=8'h4B; mem['hE3AD]=8'h0D; mem['hE3AE]=8'h00; mem['hE3AF]=8'h0D;
    mem['hE3B0]=8'h42; mem['hE3B1]=8'h52; mem['hE3B2]=8'h45; mem['hE3B3]=8'h41;
    mem['hE3B4]=8'h4B; mem['hE3B5]=8'h00; mem['hE3B6]=8'h30; mem['hE3B7]=8'h64;
    mem['hE3B8]=8'hC6; mem['hE3B9]=8'h12; mem['hE3BA]=8'h9F; mem['hE3BB]=8'h0F;
    mem['hE3BC]=8'hA6; mem['hE3BD]=8'h84; mem['hE3BE]=8'h80; mem['hE3BF]=8'h80;
    mem['hE3C0]=8'h26; mem['hE3C1]=8'h15; mem['hE3C2]=8'hAE; mem['hE3C3]=8'h01;
    mem['hE3C4]=8'h9F; mem['hE3C5]=8'h11; mem['hE3C6]=8'h9E; mem['hE3C7]=8'h3B;
    mem['hE3C8]=8'h27; mem['hE3C9]=8'h09; mem['hE3CA]=8'h9C; mem['hE3CB]=8'h11;
    mem['hE3CC]=8'h27; mem['hE3CD]=8'h09; mem['hE3CE]=8'h9E; mem['hE3CF]=8'h0F;
    mem['hE3D0]=8'h3A; mem['hE3D1]=8'h20; mem['hE3D2]=8'hE5; mem['hE3D3]=8'h9E;
    mem['hE3D4]=8'h11; mem['hE3D5]=8'h9F; mem['hE3D6]=8'h3B; mem['hE3D7]=8'h9E;
    mem['hE3D8]=8'h0F; mem['hE3D9]=8'h4D; mem['hE3DA]=8'h39; mem['hE3DB]=8'h8D;
    mem['hE3DC]=8'h17; mem['hE3DD]=8'hDE; mem['hE3DE]=8'h41; mem['hE3DF]=8'h33;
    mem['hE3E0]=8'h41; mem['hE3E1]=8'h9E; mem['hE3E2]=8'h43; mem['hE3E3]=8'h30;
    mem['hE3E4]=8'h01; mem['hE3E5]=8'hA6; mem['hE3E6]=8'h82; mem['hE3E7]=8'h36;
    mem['hE3E8]=8'h02; mem['hE3E9]=8'h9C; mem['hE3EA]=8'h47; mem['hE3EB]=8'h26;
    mem['hE3EC]=8'hF8; mem['hE3ED]=8'hDF; mem['hE3EE]=8'h45; mem['hE3EF]=8'h39;
    mem['hE3F0]=8'h4F; mem['hE3F1]=8'h58; mem['hE3F2]=8'hD3; mem['hE3F3]=8'h1F;
    mem['hE3F4]=8'hC3; mem['hE3F5]=8'h00; mem['hE3F6]=8'h3A; mem['hE3F7]=8'h25;
    mem['hE3F8]=8'h08; mem['hE3F9]=8'h10; mem['hE3FA]=8'hDF; mem['hE3FB]=8'h17;
    mem['hE3FC]=8'h10; mem['hE3FD]=8'h93; mem['hE3FE]=8'h17; mem['hE3FF]=8'h25;
    mem['hE400]=8'hEE; mem['hE401]=8'hC6; mem['hE402]=8'h0C; mem['hE403]=8'hBD;
    mem['hE404]=8'hE4; mem['hE405]=8'hD4; mem['hE406]=8'hBD; mem['hE407]=8'hF0;
    mem['hE408]=8'hA6; mem['hE409]=8'hBD; mem['hE40A]=8'hF0; mem['hE40B]=8'hF5;
    mem['hE40C]=8'h8E; mem['hE40D]=8'hE3; mem['hE40E]=8'h68; mem['hE40F]=8'h3A;
    mem['hE410]=8'h8D; mem['hE411]=8'h31; mem['hE412]=8'h8D; mem['hE413]=8'h2F;
    mem['hE414]=8'h8E; mem['hE415]=8'hE3; mem['hE416]=8'h9D; mem['hE417]=8'hBD;
    mem['hE418]=8'hF0; mem['hE419]=8'hE2; mem['hE41A]=8'h96; mem['hE41B]=8'h68;
    mem['hE41C]=8'h4C; mem['hE41D]=8'h27; mem['hE41E]=8'h03; mem['hE41F]=8'hBD;
    mem['hE420]=8'hF5; mem['hE421]=8'h0B; mem['hE422]=8'hBD; mem['hE423]=8'hF0;
    mem['hE424]=8'hA6; mem['hE425]=8'h8E; mem['hE426]=8'hE3; mem['hE427]=8'hAA;
    mem['hE428]=8'hBD; mem['hE429]=8'hF0; mem['hE42A]=8'hE2; mem['hE42B]=8'hBD;
    mem['hE42C]=8'hE1; mem['hE42D]=8'h3E; mem['hE42E]=8'hCE; mem['hE42F]=8'hFF;
    mem['hE430]=8'hFF; mem['hE431]=8'hDF; mem['hE432]=8'h68; mem['hE433]=8'h25;
    mem['hE434]=8'hF6; mem['hE435]=8'h9F; mem['hE436]=8'h83; mem['hE437]=8'h9D;
    mem['hE438]=8'h7C; mem['hE439]=8'h27; mem['hE43A]=8'hF0; mem['hE43B]=8'h25;
    mem['hE43C]=8'h0B; mem['hE43D]=8'hBD; mem['hE43E]=8'hEF; mem['hE43F]=8'h97;
    mem['hE440]=8'h7E; mem['hE441]=8'hE5; mem['hE442]=8'h71; mem['hE443]=8'hA6;
    mem['hE444]=8'h80; mem['hE445]=8'h7E; mem['hE446]=8'hF0; mem['hE447]=8'hF7;
    mem['hE448]=8'hBD; mem['hE449]=8'hE7; mem['hE44A]=8'h14; mem['hE44B]=8'h9E;
    mem['hE44C]=8'h2B; mem['hE44D]=8'h9F; mem['hE44E]=8'hF1; mem['hE44F]=8'hBD;
    mem['hE450]=8'hEF; mem['hE451]=8'h97; mem['hE452]=8'hD7; mem['hE453]=8'h03;
    mem['hE454]=8'h8D; mem['hE455]=8'h4C; mem['hE456]=8'h25; mem['hE457]=8'h12;
    mem['hE458]=8'hDC; mem['hE459]=8'h47; mem['hE45A]=8'hA3; mem['hE45B]=8'h84;
    mem['hE45C]=8'hD3; mem['hE45D]=8'h1B; mem['hE45E]=8'hDD; mem['hE45F]=8'h1B;
    mem['hE460]=8'hEE; mem['hE461]=8'h84; mem['hE462]=8'h37; mem['hE463]=8'h02;
    mem['hE464]=8'hA7; mem['hE465]=8'h80; mem['hE466]=8'h9C; mem['hE467]=8'h1B;
    mem['hE468]=8'h26; mem['hE469]=8'hF8; mem['hE46A]=8'h96; mem['hE46B]=8'hF3;
    mem['hE46C]=8'h27; mem['hE46D]=8'h1C; mem['hE46E]=8'hDC; mem['hE46F]=8'h1B;
    mem['hE470]=8'hDD; mem['hE471]=8'h43; mem['hE472]=8'hDB; mem['hE473]=8'h03;
    mem['hE474]=8'h89; mem['hE475]=8'h00; mem['hE476]=8'hDD; mem['hE477]=8'h41;
    mem['hE478]=8'hBD; mem['hE479]=8'hE3; mem['hE47A]=8'hDB; mem['hE47B]=8'hCE;
    mem['hE47C]=8'h00; mem['hE47D]=8'hEF; mem['hE47E]=8'h37; mem['hE47F]=8'h02;
    mem['hE480]=8'hA7; mem['hE481]=8'h80; mem['hE482]=8'h9C; mem['hE483]=8'h45;
    mem['hE484]=8'h26; mem['hE485]=8'hF8; mem['hE486]=8'h9E; mem['hE487]=8'h41;
    mem['hE488]=8'h9F; mem['hE489]=8'h1B; mem['hE48A]=8'h8D; mem['hE48B]=8'h36;
    mem['hE48C]=8'h8D; mem['hE48D]=8'h02; mem['hE48E]=8'h20; mem['hE48F]=8'h9B;
    mem['hE490]=8'h9E; mem['hE491]=8'h19; mem['hE492]=8'hEC; mem['hE493]=8'h84;
    mem['hE494]=8'h27; mem['hE495]=8'h21; mem['hE496]=8'h33; mem['hE497]=8'h04;
    mem['hE498]=8'hA6; mem['hE499]=8'hC0; mem['hE49A]=8'h26; mem['hE49B]=8'hFC;
    mem['hE49C]=8'hEF; mem['hE49D]=8'h84; mem['hE49E]=8'hAE; mem['hE49F]=8'h84;
    mem['hE4A0]=8'h20; mem['hE4A1]=8'hF0; mem['hE4A2]=8'hDC; mem['hE4A3]=8'h2B;
    mem['hE4A4]=8'h9E; mem['hE4A5]=8'h19; mem['hE4A6]=8'hEE; mem['hE4A7]=8'h84;
    mem['hE4A8]=8'h27; mem['hE4A9]=8'h09; mem['hE4AA]=8'h10; mem['hE4AB]=8'hA3;
    mem['hE4AC]=8'h02; mem['hE4AD]=8'h23; mem['hE4AE]=8'h06; mem['hE4AF]=8'hAE;
    mem['hE4B0]=8'h84; mem['hE4B1]=8'h20; mem['hE4B2]=8'hF3; mem['hE4B3]=8'h1A;
    mem['hE4B4]=8'h01; mem['hE4B5]=8'h9F; mem['hE4B6]=8'h47; mem['hE4B7]=8'h39;
    mem['hE4B8]=8'h26; mem['hE4B9]=8'hFB; mem['hE4BA]=8'h9E; mem['hE4BB]=8'h19;
    mem['hE4BC]=8'h6F; mem['hE4BD]=8'h80; mem['hE4BE]=8'h6F; mem['hE4BF]=8'h80;
    mem['hE4C0]=8'h9F; mem['hE4C1]=8'h1B; mem['hE4C2]=8'h9E; mem['hE4C3]=8'h19;
    mem['hE4C4]=8'hBD; mem['hE4C5]=8'hE6; mem['hE4C6]=8'h68; mem['hE4C7]=8'h9E;
    mem['hE4C8]=8'h27; mem['hE4C9]=8'h9F; mem['hE4CA]=8'h23; mem['hE4CB]=8'hBD;
    mem['hE4CC]=8'hE5; mem['hE4CD]=8'h9C; mem['hE4CE]=8'h9E; mem['hE4CF]=8'h1B;
    mem['hE4D0]=8'h9F; mem['hE4D1]=8'h1D; mem['hE4D2]=8'h9F; mem['hE4D3]=8'h1F;
    mem['hE4D4]=8'h8E; mem['hE4D5]=8'h00; mem['hE4D6]=8'hC9; mem['hE4D7]=8'h9F;
    mem['hE4D8]=8'h0B; mem['hE4D9]=8'hAE; mem['hE4DA]=8'hE4; mem['hE4DB]=8'h10;
    mem['hE4DC]=8'hDE; mem['hE4DD]=8'h21; mem['hE4DE]=8'h6F; mem['hE4DF]=8'hE2;
    mem['hE4E0]=8'h0F; mem['hE4E1]=8'h2D; mem['hE4E2]=8'h0F; mem['hE4E3]=8'h2E;
    mem['hE4E4]=8'h0F; mem['hE4E5]=8'h08; mem['hE4E6]=8'h6E; mem['hE4E7]=8'h84;
    mem['hE4E8]=8'h86; mem['hE4E9]=8'h80; mem['hE4EA]=8'h97; mem['hE4EB]=8'h08;
    mem['hE4EC]=8'hBD; mem['hE4ED]=8'hE7; mem['hE4EE]=8'h36; mem['hE4EF]=8'hBD;
    mem['hE4F0]=8'hE3; mem['hE4F1]=8'hB6; mem['hE4F2]=8'h32; mem['hE4F3]=8'h62;
    mem['hE4F4]=8'h26; mem['hE4F5]=8'h04; mem['hE4F6]=8'h9E; mem['hE4F7]=8'h0F;
    mem['hE4F8]=8'h32; mem['hE4F9]=8'h85; mem['hE4FA]=8'hC6; mem['hE4FB]=8'h09;
    mem['hE4FC]=8'hBD; mem['hE4FD]=8'hE3; mem['hE4FE]=8'hF0; mem['hE4FF]=8'hBD;
    mem['hE500]=8'hE6; mem['hE501]=8'h95; mem['hE502]=8'hDC; mem['hE503]=8'h68;
    mem['hE504]=8'h34; mem['hE505]=8'h16; mem['hE506]=8'hC6; mem['hE507]=8'hA0;
    mem['hE508]=8'hBD; mem['hE509]=8'hE9; mem['hE50A]=8'hF8; mem['hE50B]=8'hBD;
    mem['hE50C]=8'hE8; mem['hE50D]=8'hCC; mem['hE50E]=8'hBD; mem['hE50F]=8'hE8;
    mem['hE510]=8'hCA; mem['hE511]=8'hD6; mem['hE512]=8'h54; mem['hE513]=8'hCA;
    mem['hE514]=8'h7F; mem['hE515]=8'hD4; mem['hE516]=8'h50; mem['hE517]=8'hD7;
    mem['hE518]=8'h50; mem['hE519]=8'h10; mem['hE51A]=8'h8E; mem['hE51B]=8'hE5;
    mem['hE51C]=8'h20; mem['hE51D]=8'h7E; mem['hE51E]=8'hE9; mem['hE51F]=8'h73;
    mem['hE520]=8'h8E; mem['hE521]=8'hF2; mem['hE522]=8'h0B; mem['hE523]=8'hBD;
    mem['hE524]=8'hF3; mem['hE525]=8'h5A; mem['hE526]=8'h9D; mem['hE527]=8'h82;
    mem['hE528]=8'h81; mem['hE529]=8'hA4; mem['hE52A]=8'h26; mem['hE52B]=8'h05;
    mem['hE52C]=8'h9D; mem['hE52D]=8'h7C; mem['hE52E]=8'hBD; mem['hE52F]=8'hE8;
    mem['hE530]=8'hCA; mem['hE531]=8'hBD; mem['hE532]=8'hF3; mem['hE533]=8'hB3;
    mem['hE534]=8'hBD; mem['hE535]=8'hE9; mem['hE536]=8'h6F; mem['hE537]=8'hDC;
    mem['hE538]=8'h3B; mem['hE539]=8'h34; mem['hE53A]=8'h06; mem['hE53B]=8'h86;
    mem['hE53C]=8'h80; mem['hE53D]=8'h34; mem['hE53E]=8'h02; mem['hE53F]=8'h1C;
    mem['hE540]=8'hAF; mem['hE541]=8'h8D; mem['hE542]=8'h60; mem['hE543]=8'h9E;
    mem['hE544]=8'h83; mem['hE545]=8'h9F; mem['hE546]=8'h2F; mem['hE547]=8'hA6;
    mem['hE548]=8'h80; mem['hE549]=8'h27; mem['hE54A]=8'h07; mem['hE54B]=8'h81;
    mem['hE54C]=8'h3A; mem['hE54D]=8'h27; mem['hE54E]=8'h22; mem['hE54F]=8'h7E;
    mem['hE550]=8'hEA; mem['hE551]=8'h00; mem['hE552]=8'hA6; mem['hE553]=8'h81;
    mem['hE554]=8'h97; mem['hE555]=8'h00; mem['hE556]=8'h27; mem['hE557]=8'h72;
    mem['hE558]=8'hEC; mem['hE559]=8'h80; mem['hE55A]=8'hDD; mem['hE55B]=8'h68;
    mem['hE55C]=8'h9F; mem['hE55D]=8'h83; mem['hE55E]=8'h96; mem['hE55F]=8'h8C;
    mem['hE560]=8'h27; mem['hE561]=8'h0F; mem['hE562]=8'h86; mem['hE563]=8'h5B;
    mem['hE564]=8'hBD; mem['hE565]=8'hE0; mem['hE566]=8'h14; mem['hE567]=8'h96;
    mem['hE568]=8'h68; mem['hE569]=8'hBD; mem['hE56A]=8'hF5; mem['hE56B]=8'h12;
    mem['hE56C]=8'h86; mem['hE56D]=8'h5D; mem['hE56E]=8'hBD; mem['hE56F]=8'hE0;
    mem['hE570]=8'h14; mem['hE571]=8'h9D; mem['hE572]=8'h7C; mem['hE573]=8'h8D;
    mem['hE574]=8'h02; mem['hE575]=8'h20; mem['hE576]=8'hC8; mem['hE577]=8'h27;
    mem['hE578]=8'h29; mem['hE579]=8'h4D; mem['hE57A]=8'h10; mem['hE57B]=8'h2A;
    mem['hE57C]=8'h01; mem['hE57D]=8'hB8; mem['hE57E]=8'h81; mem['hE57F]=8'hFF;
    mem['hE580]=8'h27; mem['hE581]=8'h0F; mem['hE582]=8'h81; mem['hE583]=8'h9E;
    mem['hE584]=8'h22; mem['hE585]=8'hC9; mem['hE586]=8'hBE; mem['hE587]=8'hE0;
    mem['hE588]=8'hF1; mem['hE589]=8'h48; mem['hE58A]=8'h1F; mem['hE58B]=8'h89;
    mem['hE58C]=8'h3A; mem['hE58D]=8'h9D; mem['hE58E]=8'h7C; mem['hE58F]=8'h6E;
    mem['hE590]=8'h94; mem['hE591]=8'h9D; mem['hE592]=8'h7C; mem['hE593]=8'h81;
    mem['hE594]=8'h97; mem['hE595]=8'h10; mem['hE596]=8'h27; mem['hE597]=8'h14;
    mem['hE598]=8'hED; mem['hE599]=8'h7E; mem['hE59A]=8'hEA; mem['hE59B]=8'h00;
    mem['hE59C]=8'h9E; mem['hE59D]=8'h19; mem['hE59E]=8'h30; mem['hE59F]=8'h1F;
    mem['hE5A0]=8'h9F; mem['hE5A1]=8'h33; mem['hE5A2]=8'h39; mem['hE5A3]=8'hBD;
    mem['hE5A4]=8'hE0; mem['hE5A5]=8'h05; mem['hE5A6]=8'h27; mem['hE5A7]=8'h0A;
    mem['hE5A8]=8'h81; mem['hE5A9]=8'h03; mem['hE5AA]=8'h27; mem['hE5AB]=8'h12;
    mem['hE5AC]=8'h81; mem['hE5AD]=8'h13; mem['hE5AE]=8'h27; mem['hE5AF]=8'h03;
    mem['hE5B0]=8'h97; mem['hE5B1]=8'h73; mem['hE5B2]=8'h39; mem['hE5B3]=8'hBD;
    mem['hE5B4]=8'hE0; mem['hE5B5]=8'h05; mem['hE5B6]=8'h27; mem['hE5B7]=8'hFB;
    mem['hE5B8]=8'h20; mem['hE5B9]=8'hEE; mem['hE5BA]=8'h9D; mem['hE5BB]=8'h82;
    mem['hE5BC]=8'h20; mem['hE5BD]=8'h02; mem['hE5BE]=8'h1A; mem['hE5BF]=8'h01;
    mem['hE5C0]=8'h26; mem['hE5C1]=8'h31; mem['hE5C2]=8'h9E; mem['hE5C3]=8'h83;
    mem['hE5C4]=8'h9F; mem['hE5C5]=8'h2F; mem['hE5C6]=8'h06; mem['hE5C7]=8'h00;
    mem['hE5C8]=8'h32; mem['hE5C9]=8'h62; mem['hE5CA]=8'h9E; mem['hE5CB]=8'h68;
    mem['hE5CC]=8'h8C; mem['hE5CD]=8'hFF; mem['hE5CE]=8'hFF; mem['hE5CF]=8'h27;
    mem['hE5D0]=8'h06; mem['hE5D1]=8'h9F; mem['hE5D2]=8'h29; mem['hE5D3]=8'h9E;
    mem['hE5D4]=8'h2F; mem['hE5D5]=8'h9F; mem['hE5D6]=8'h2D; mem['hE5D7]=8'h8E;
    mem['hE5D8]=8'hE3; mem['hE5D9]=8'hAE; mem['hE5DA]=8'h0D; mem['hE5DB]=8'h00;
    mem['hE5DC]=8'h10; mem['hE5DD]=8'h2A; mem['hE5DE]=8'hFE; mem['hE5DF]=8'h42;
    mem['hE5E0]=8'h7E; mem['hE5E1]=8'hE4; mem['hE5E2]=8'h17; mem['hE5E3]=8'h26;
    mem['hE5E4]=8'h0E; mem['hE5E5]=8'hC6; mem['hE5E6]=8'h20; mem['hE5E7]=8'h9E;
    mem['hE5E8]=8'h2D; mem['hE5E9]=8'h10; mem['hE5EA]=8'h27; mem['hE5EB]=8'hFE;
    mem['hE5EC]=8'h16; mem['hE5ED]=8'h9F; mem['hE5EE]=8'h83; mem['hE5EF]=8'h9E;
    mem['hE5F0]=8'h29; mem['hE5F1]=8'h9F; mem['hE5F2]=8'h68; mem['hE5F3]=8'h39;
    mem['hE5F4]=8'h27; mem['hE5F5]=8'h2C; mem['hE5F6]=8'hBD; mem['hE5F7]=8'hEB;
    mem['hE5F8]=8'h6A; mem['hE5F9]=8'h34; mem['hE5FA]=8'h06; mem['hE5FB]=8'h9E;
    mem['hE5FC]=8'h27; mem['hE5FD]=8'h9D; mem['hE5FE]=8'h82; mem['hE5FF]=8'h27;
    mem['hE600]=8'h0C; mem['hE601]=8'hBD; mem['hE602]=8'hE9; mem['hE603]=8'hF6;
    mem['hE604]=8'hBD; mem['hE605]=8'hEE; mem['hE606]=8'hC1; mem['hE607]=8'h30;
    mem['hE608]=8'h1F; mem['hE609]=8'h9C; mem['hE60A]=8'h71; mem['hE60B]=8'h22;
    mem['hE60C]=8'h18; mem['hE60D]=8'h1F; mem['hE60E]=8'h10; mem['hE60F]=8'hA3;
    mem['hE610]=8'hE1; mem['hE611]=8'h25; mem['hE612]=8'h12; mem['hE613]=8'h1F;
    mem['hE614]=8'h03; mem['hE615]=8'h83; mem['hE616]=8'h00; mem['hE617]=8'h3A;
    mem['hE618]=8'h25; mem['hE619]=8'h0B; mem['hE61A]=8'h93; mem['hE61B]=8'h1B;
    mem['hE61C]=8'h25; mem['hE61D]=8'h07; mem['hE61E]=8'hDF; mem['hE61F]=8'h21;
    mem['hE620]=8'h9F; mem['hE621]=8'h27; mem['hE622]=8'h7E; mem['hE623]=8'hE4;
    mem['hE624]=8'hC7; mem['hE625]=8'h7E; mem['hE626]=8'hE4; mem['hE627]=8'h01;
    mem['hE628]=8'h9D; mem['hE629]=8'h82; mem['hE62A]=8'h10; mem['hE62B]=8'h27;
    mem['hE62C]=8'hFE; mem['hE62D]=8'h94; mem['hE62E]=8'hBD; mem['hE62F]=8'hE4;
    mem['hE630]=8'hC7; mem['hE631]=8'h20; mem['hE632]=8'h19; mem['hE633]=8'h1F;
    mem['hE634]=8'h89; mem['hE635]=8'h9D; mem['hE636]=8'h7C; mem['hE637]=8'hC1;
    mem['hE638]=8'hA0; mem['hE639]=8'h27; mem['hE63A]=8'h16; mem['hE63B]=8'hC1;
    mem['hE63C]=8'hA1; mem['hE63D]=8'h26; mem['hE63E]=8'h45; mem['hE63F]=8'hC6;
    mem['hE640]=8'h03; mem['hE641]=8'hBD; mem['hE642]=8'hE3; mem['hE643]=8'hF0;
    mem['hE644]=8'hDE; mem['hE645]=8'h83; mem['hE646]=8'h9E; mem['hE647]=8'h68;
    mem['hE648]=8'h86; mem['hE649]=8'hA1; mem['hE64A]=8'h34; mem['hE64B]=8'h52;
    mem['hE64C]=8'h8D; mem['hE64D]=8'h03; mem['hE64E]=8'h7E; mem['hE64F]=8'hE5;
    mem['hE650]=8'h3F; mem['hE651]=8'h9D; mem['hE652]=8'h82; mem['hE653]=8'hBD;
    mem['hE654]=8'hE7; mem['hE655]=8'h14; mem['hE656]=8'h8D; mem['hE657]=8'h40;
    mem['hE658]=8'h30; mem['hE659]=8'h01; mem['hE65A]=8'hDC; mem['hE65B]=8'h2B;
    mem['hE65C]=8'h10; mem['hE65D]=8'h93; mem['hE65E]=8'h68; mem['hE65F]=8'h22;
    mem['hE660]=8'h02; mem['hE661]=8'h9E; mem['hE662]=8'h19; mem['hE663]=8'hBD;
    mem['hE664]=8'hE4; mem['hE665]=8'hA6; mem['hE666]=8'h25; mem['hE667]=8'h17;
    mem['hE668]=8'h30; mem['hE669]=8'h1F; mem['hE66A]=8'h9F; mem['hE66B]=8'h83;
    mem['hE66C]=8'h39; mem['hE66D]=8'h26; mem['hE66E]=8'hFD; mem['hE66F]=8'h86;
    mem['hE670]=8'hFF; mem['hE671]=8'h97; mem['hE672]=8'h3B; mem['hE673]=8'hBD;
    mem['hE674]=8'hE3; mem['hE675]=8'hB6; mem['hE676]=8'h1F; mem['hE677]=8'h14;
    mem['hE678]=8'h81; mem['hE679]=8'h21; mem['hE67A]=8'h27; mem['hE67B]=8'h0B;
    mem['hE67C]=8'hC6; mem['hE67D]=8'h04; mem['hE67E]=8'h8C; mem['hE67F]=8'hC6;
    mem['hE680]=8'h0E; mem['hE681]=8'h7E; mem['hE682]=8'hE4; mem['hE683]=8'h03;
    mem['hE684]=8'h7E; mem['hE685]=8'hEA; mem['hE686]=8'h00; mem['hE687]=8'h35;
    mem['hE688]=8'h52; mem['hE689]=8'h9F; mem['hE68A]=8'h68; mem['hE68B]=8'hDF;
    mem['hE68C]=8'h83; mem['hE68D]=8'h8D; mem['hE68E]=8'h06; mem['hE68F]=8'h8C;
    mem['hE690]=8'h8D; mem['hE691]=8'h06; mem['hE692]=8'h9F; mem['hE693]=8'h83;
    mem['hE694]=8'h39; mem['hE695]=8'hC6; mem['hE696]=8'h3A; mem['hE697]=8'h86;
    mem['hE698]=8'h5F; mem['hE699]=8'hD7; mem['hE69A]=8'h01; mem['hE69B]=8'h5F;
    mem['hE69C]=8'h9E; mem['hE69D]=8'h83; mem['hE69E]=8'h1F; mem['hE69F]=8'h98;
    mem['hE6A0]=8'hD6; mem['hE6A1]=8'h01; mem['hE6A2]=8'h97; mem['hE6A3]=8'h01;
    mem['hE6A4]=8'hA6; mem['hE6A5]=8'h84; mem['hE6A6]=8'h27; mem['hE6A7]=8'hEC;
    mem['hE6A8]=8'h34; mem['hE6A9]=8'h04; mem['hE6AA]=8'hA1; mem['hE6AB]=8'hE0;
    mem['hE6AC]=8'h27; mem['hE6AD]=8'hE6; mem['hE6AE]=8'h30; mem['hE6AF]=8'h01;
    mem['hE6B0]=8'h81; mem['hE6B1]=8'h22; mem['hE6B2]=8'h27; mem['hE6B3]=8'hEA;
    mem['hE6B4]=8'h4C; mem['hE6B5]=8'h26; mem['hE6B6]=8'h02; mem['hE6B7]=8'h30;
    mem['hE6B8]=8'h01; mem['hE6B9]=8'h81; mem['hE6BA]=8'h86; mem['hE6BB]=8'h26;
    mem['hE6BC]=8'hE7; mem['hE6BD]=8'h0C; mem['hE6BE]=8'h04; mem['hE6BF]=8'h20;
    mem['hE6C0]=8'hE3; mem['hE6C1]=8'hBD; mem['hE6C2]=8'hE8; mem['hE6C3]=8'hCA;
    mem['hE6C4]=8'h9D; mem['hE6C5]=8'h82; mem['hE6C6]=8'h81; mem['hE6C7]=8'h81;
    mem['hE6C8]=8'h27; mem['hE6C9]=8'h05; mem['hE6CA]=8'hC6; mem['hE6CB]=8'hA2;
    mem['hE6CC]=8'hBD; mem['hE6CD]=8'hE9; mem['hE6CE]=8'hF8; mem['hE6CF]=8'h96;
    mem['hE6D0]=8'h4F; mem['hE6D1]=8'h26; mem['hE6D2]=8'h13; mem['hE6D3]=8'h0F;
    mem['hE6D4]=8'h04; mem['hE6D5]=8'h8D; mem['hE6D6]=8'hB6; mem['hE6D7]=8'h4D;
    mem['hE6D8]=8'h27; mem['hE6D9]=8'hBA; mem['hE6DA]=8'h9D; mem['hE6DB]=8'h7C;
    mem['hE6DC]=8'h81; mem['hE6DD]=8'h84; mem['hE6DE]=8'h26; mem['hE6DF]=8'hF5;
    mem['hE6E0]=8'h0A; mem['hE6E1]=8'h04; mem['hE6E2]=8'h2A; mem['hE6E3]=8'hF1;
    mem['hE6E4]=8'h9D; mem['hE6E5]=8'h7C; mem['hE6E6]=8'h9D; mem['hE6E7]=8'h82;
    mem['hE6E8]=8'h10; mem['hE6E9]=8'h25; mem['hE6EA]=8'hFF; mem['hE6EB]=8'h65;
    mem['hE6EC]=8'h7E; mem['hE6ED]=8'hE5; mem['hE6EE]=8'h77; mem['hE6EF]=8'hBD;
    mem['hE6F0]=8'hEE; mem['hE6F1]=8'h8F; mem['hE6F2]=8'hC6; mem['hE6F3]=8'h81;
    mem['hE6F4]=8'hBD; mem['hE6F5]=8'hE9; mem['hE6F6]=8'hF8; mem['hE6F7]=8'h34;
    mem['hE6F8]=8'h02; mem['hE6F9]=8'h81; mem['hE6FA]=8'hA1; mem['hE6FB]=8'h27;
    mem['hE6FC]=8'h04; mem['hE6FD]=8'h81; mem['hE6FE]=8'hA0; mem['hE6FF]=8'h26;
    mem['hE700]=8'h83; mem['hE701]=8'h0A; mem['hE702]=8'h53; mem['hE703]=8'h26;
    mem['hE704]=8'h05; mem['hE705]=8'h35; mem['hE706]=8'h04; mem['hE707]=8'h7E;
    mem['hE708]=8'hE6; mem['hE709]=8'h35; mem['hE70A]=8'h9D; mem['hE70B]=8'h7C;
    mem['hE70C]=8'h8D; mem['hE70D]=8'h06; mem['hE70E]=8'h81; mem['hE70F]=8'h2C;
    mem['hE710]=8'h27; mem['hE711]=8'hEF; mem['hE712]=8'h35; mem['hE713]=8'h84;
    mem['hE714]=8'h9E; mem['hE715]=8'h74; mem['hE716]=8'h9F; mem['hE717]=8'h2B;
    mem['hE718]=8'h24; mem['hE719]=8'h61; mem['hE71A]=8'h80; mem['hE71B]=8'h30;
    mem['hE71C]=8'h97; mem['hE71D]=8'h01; mem['hE71E]=8'hDC; mem['hE71F]=8'h2B;
    mem['hE720]=8'h81; mem['hE721]=8'h18; mem['hE722]=8'h22; mem['hE723]=8'hDB;
    mem['hE724]=8'h58; mem['hE725]=8'h49; mem['hE726]=8'h58; mem['hE727]=8'h49;
    mem['hE728]=8'hD3; mem['hE729]=8'h2B; mem['hE72A]=8'h58; mem['hE72B]=8'h49;
    mem['hE72C]=8'hDB; mem['hE72D]=8'h01; mem['hE72E]=8'h89; mem['hE72F]=8'h00;
    mem['hE730]=8'hDD; mem['hE731]=8'h2B; mem['hE732]=8'h9D; mem['hE733]=8'h7C;
    mem['hE734]=8'h20; mem['hE735]=8'hE2; mem['hE736]=8'hBD; mem['hE737]=8'hEA;
    mem['hE738]=8'hDB; mem['hE739]=8'h9F; mem['hE73A]=8'h3B; mem['hE73B]=8'hC6;
    mem['hE73C]=8'hAE; mem['hE73D]=8'hBD; mem['hE73E]=8'hE9; mem['hE73F]=8'hF8;
    mem['hE740]=8'h96; mem['hE741]=8'h06; mem['hE742]=8'h34; mem['hE743]=8'h02;
    mem['hE744]=8'hBD; mem['hE745]=8'hE8; mem['hE746]=8'hDF; mem['hE747]=8'h35;
    mem['hE748]=8'h02; mem['hE749]=8'h46; mem['hE74A]=8'hBD; mem['hE74B]=8'hE8;
    mem['hE74C]=8'hD1; mem['hE74D]=8'h10; mem['hE74E]=8'h27; mem['hE74F]=8'h0C;
    mem['hE750]=8'h28; mem['hE751]=8'h9E; mem['hE752]=8'h52; mem['hE753]=8'hDC;
    mem['hE754]=8'h21; mem['hE755]=8'h10; mem['hE756]=8'hA3; mem['hE757]=8'h02;
    mem['hE758]=8'h24; mem['hE759]=8'h11; mem['hE75A]=8'h9C; mem['hE75B]=8'h1B;
    mem['hE75C]=8'h25; mem['hE75D]=8'h0D; mem['hE75E]=8'hE6; mem['hE75F]=8'h84;
    mem['hE760]=8'hBD; mem['hE761]=8'hEC; mem['hE762]=8'h91; mem['hE763]=8'h9E;
    mem['hE764]=8'h4D; mem['hE765]=8'hBD; mem['hE766]=8'hED; mem['hE767]=8'hC7;
    mem['hE768]=8'h8E; mem['hE769]=8'h00; mem['hE76A]=8'h56; mem['hE76B]=8'h9F;
    mem['hE76C]=8'h4D; mem['hE76D]=8'hBD; mem['hE76E]=8'hED; mem['hE76F]=8'hF9;
    mem['hE770]=8'hDE; mem['hE771]=8'h4D; mem['hE772]=8'h9E; mem['hE773]=8'h3B;
    mem['hE774]=8'h37; mem['hE775]=8'h26; mem['hE776]=8'hA7; mem['hE777]=8'h84;
    mem['hE778]=8'h10; mem['hE779]=8'hAF; mem['hE77A]=8'h02; mem['hE77B]=8'h39;
    mem['hE77C]=8'h3F; mem['hE77D]=8'h52; mem['hE77E]=8'h45; mem['hE77F]=8'h44;
    mem['hE780]=8'h4F; mem['hE781]=8'h0D; mem['hE782]=8'h00; mem['hE783]=8'h7E;
    mem['hE784]=8'hE4; mem['hE785]=8'h03; mem['hE786]=8'h96; mem['hE787]=8'h09;
    mem['hE788]=8'h27; mem['hE789]=8'h07; mem['hE78A]=8'h9E; mem['hE78B]=8'h31;
    mem['hE78C]=8'h9F; mem['hE78D]=8'h68; mem['hE78E]=8'h7E; mem['hE78F]=8'hEA;
    mem['hE790]=8'h00; mem['hE791]=8'h8E; mem['hE792]=8'hE7; mem['hE793]=8'h7B;
    mem['hE794]=8'hBD; mem['hE795]=8'hF0; mem['hE796]=8'hE2; mem['hE797]=8'h9E;
    mem['hE798]=8'h2F; mem['hE799]=8'h9F; mem['hE79A]=8'h83; mem['hE79B]=8'h39;
    mem['hE79C]=8'hC6; mem['hE79D]=8'h16; mem['hE79E]=8'h9E; mem['hE79F]=8'h68;
    mem['hE7A0]=8'h30; mem['hE7A1]=8'h01; mem['hE7A2]=8'h27; mem['hE7A3]=8'hDF;
    mem['hE7A4]=8'h8D; mem['hE7A5]=8'h01; mem['hE7A6]=8'h39; mem['hE7A7]=8'h81;
    mem['hE7A8]=8'h22; mem['hE7A9]=8'h26; mem['hE7AA]=8'h0B; mem['hE7AB]=8'hBD;
    mem['hE7AC]=8'hE9; mem['hE7AD]=8'hCD; mem['hE7AE]=8'hC6; mem['hE7AF]=8'h3B;
    mem['hE7B0]=8'hBD; mem['hE7B1]=8'hE9; mem['hE7B2]=8'hF8; mem['hE7B3]=8'hBD;
    mem['hE7B4]=8'hF0; mem['hE7B5]=8'hE5; mem['hE7B6]=8'h8E; mem['hE7B7]=8'h00;
    mem['hE7B8]=8'hF3; mem['hE7B9]=8'h6F; mem['hE7BA]=8'h84; mem['hE7BB]=8'h8D;
    mem['hE7BC]=8'h06; mem['hE7BD]=8'hC6; mem['hE7BE]=8'h2C; mem['hE7BF]=8'hE7;
    mem['hE7C0]=8'h84; mem['hE7C1]=8'h20; mem['hE7C2]=8'h16; mem['hE7C3]=8'hBD;
    mem['hE7C4]=8'hF0; mem['hE7C5]=8'hF5; mem['hE7C6]=8'hBD; mem['hE7C7]=8'hF0;
    mem['hE7C8]=8'hF2; mem['hE7C9]=8'hBD; mem['hE7CA]=8'hE1; mem['hE7CB]=8'h3E;
    mem['hE7CC]=8'h24; mem['hE7CD]=8'h05; mem['hE7CE]=8'h32; mem['hE7CF]=8'h64;
    mem['hE7D0]=8'h7E; mem['hE7D1]=8'hE5; mem['hE7D2]=8'hC6; mem['hE7D3]=8'hC6;
    mem['hE7D4]=8'h2E; mem['hE7D5]=8'h39; mem['hE7D6]=8'h9E; mem['hE7D7]=8'h33;
    mem['hE7D8]=8'h86; mem['hE7D9]=8'h4F; mem['hE7DA]=8'h97; mem['hE7DB]=8'h09;
    mem['hE7DC]=8'h9F; mem['hE7DD]=8'h35; mem['hE7DE]=8'hBD; mem['hE7DF]=8'hEA;
    mem['hE7E0]=8'hDB; mem['hE7E1]=8'h9F; mem['hE7E2]=8'h3B; mem['hE7E3]=8'h9E;
    mem['hE7E4]=8'h83; mem['hE7E5]=8'h9F; mem['hE7E6]=8'h2B; mem['hE7E7]=8'h9E;
    mem['hE7E8]=8'h35; mem['hE7E9]=8'hA6; mem['hE7EA]=8'h84; mem['hE7EB]=8'h26;
    mem['hE7EC]=8'h09; mem['hE7ED]=8'h96; mem['hE7EE]=8'h09; mem['hE7EF]=8'h26;
    mem['hE7F0]=8'h51; mem['hE7F1]=8'hBD; mem['hE7F2]=8'hF0; mem['hE7F3]=8'hF5;
    mem['hE7F4]=8'h8D; mem['hE7F5]=8'hCD; mem['hE7F6]=8'h9F; mem['hE7F7]=8'h83;
    mem['hE7F8]=8'h9D; mem['hE7F9]=8'h7C; mem['hE7FA]=8'hD6; mem['hE7FB]=8'h06;
    mem['hE7FC]=8'h27; mem['hE7FD]=8'h23; mem['hE7FE]=8'h9E; mem['hE7FF]=8'h83;
    mem['hE800]=8'h97; mem['hE801]=8'h01; mem['hE802]=8'h81; mem['hE803]=8'h22;
    mem['hE804]=8'h27; mem['hE805]=8'h0E; mem['hE806]=8'h30; mem['hE807]=8'h1F;
    mem['hE808]=8'h4F; mem['hE809]=8'h97; mem['hE80A]=8'h01; mem['hE80B]=8'hBD;
    mem['hE80C]=8'hE1; mem['hE80D]=8'h30; mem['hE80E]=8'h86; mem['hE80F]=8'h3A;
    mem['hE810]=8'h97; mem['hE811]=8'h01; mem['hE812]=8'h86; mem['hE813]=8'h2C;
    mem['hE814]=8'h97; mem['hE815]=8'h02; mem['hE816]=8'hBD; mem['hE817]=8'hEC;
    mem['hE818]=8'hA2; mem['hE819]=8'hBD; mem['hE81A]=8'hE9; mem['hE81B]=8'hD2;
    mem['hE81C]=8'hBD; mem['hE81D]=8'hE7; mem['hE81E]=8'h51; mem['hE81F]=8'h20;
    mem['hE820]=8'h06; mem['hE821]=8'hBD; mem['hE822]=8'hF4; mem['hE823]=8'h58;
    mem['hE824]=8'hBD; mem['hE825]=8'hF3; mem['hE826]=8'h79; mem['hE827]=8'h9D;
    mem['hE828]=8'h82; mem['hE829]=8'h27; mem['hE82A]=8'h06; mem['hE82B]=8'h81;
    mem['hE82C]=8'h2C; mem['hE82D]=8'h10; mem['hE82E]=8'h26; mem['hE82F]=8'hFF;
    mem['hE830]=8'h52; mem['hE831]=8'h9E; mem['hE832]=8'h83; mem['hE833]=8'h9F;
    mem['hE834]=8'h35; mem['hE835]=8'h9E; mem['hE836]=8'h2B; mem['hE837]=8'h9F;
    mem['hE838]=8'h83; mem['hE839]=8'h9D; mem['hE83A]=8'h82; mem['hE83B]=8'h27;
    mem['hE83C]=8'h21; mem['hE83D]=8'hBD; mem['hE83E]=8'hE9; mem['hE83F]=8'hF6;
    mem['hE840]=8'h20; mem['hE841]=8'h9C; mem['hE842]=8'h9F; mem['hE843]=8'h83;
    mem['hE844]=8'hBD; mem['hE845]=8'hE6; mem['hE846]=8'h95; mem['hE847]=8'h30;
    mem['hE848]=8'h01; mem['hE849]=8'h4D; mem['hE84A]=8'h26; mem['hE84B]=8'h0A;
    mem['hE84C]=8'hC6; mem['hE84D]=8'h06; mem['hE84E]=8'hEE; mem['hE84F]=8'h81;
    mem['hE850]=8'h27; mem['hE851]=8'h41; mem['hE852]=8'hEC; mem['hE853]=8'h81;
    mem['hE854]=8'hDD; mem['hE855]=8'h31; mem['hE856]=8'hA6; mem['hE857]=8'h84;
    mem['hE858]=8'h81; mem['hE859]=8'h86; mem['hE85A]=8'h26; mem['hE85B]=8'hE6;
    mem['hE85C]=8'h20; mem['hE85D]=8'h98; mem['hE85E]=8'h9E; mem['hE85F]=8'h35;
    mem['hE860]=8'hD6; mem['hE861]=8'h09; mem['hE862]=8'h10; mem['hE863]=8'h26;
    mem['hE864]=8'hFD; mem['hE865]=8'h3A; mem['hE866]=8'hA6; mem['hE867]=8'h84;
    mem['hE868]=8'h27; mem['hE869]=8'h06; mem['hE86A]=8'h8E; mem['hE86B]=8'hE8;
    mem['hE86C]=8'h70; mem['hE86D]=8'h7E; mem['hE86E]=8'hF0; mem['hE86F]=8'hE2;
    mem['hE870]=8'h39; mem['hE871]=8'h3F; mem['hE872]=8'h45; mem['hE873]=8'h58;
    mem['hE874]=8'h54; mem['hE875]=8'h52; mem['hE876]=8'h41; mem['hE877]=8'h20;
    mem['hE878]=8'h49; mem['hE879]=8'h47; mem['hE87A]=8'h4E; mem['hE87B]=8'h4F;
    mem['hE87C]=8'h52; mem['hE87D]=8'h45; mem['hE87E]=8'h44; mem['hE87F]=8'h0D;
    mem['hE880]=8'h00; mem['hE881]=8'h26; mem['hE882]=8'h04; mem['hE883]=8'h9E;
    mem['hE884]=8'h74; mem['hE885]=8'h20; mem['hE886]=8'h03; mem['hE887]=8'hBD;
    mem['hE888]=8'hEA; mem['hE889]=8'hDB; mem['hE88A]=8'h9F; mem['hE88B]=8'h3B;
    mem['hE88C]=8'hBD; mem['hE88D]=8'hE3; mem['hE88E]=8'hB6; mem['hE88F]=8'h27;
    mem['hE890]=8'h04; mem['hE891]=8'hC6; mem['hE892]=8'h00; mem['hE893]=8'h20;
    mem['hE894]=8'h47; mem['hE895]=8'h1F; mem['hE896]=8'h14; mem['hE897]=8'h30;
    mem['hE898]=8'h03; mem['hE899]=8'hBD; mem['hE89A]=8'hF3; mem['hE89B]=8'h5A;
    mem['hE89C]=8'hA6; mem['hE89D]=8'h68; mem['hE89E]=8'h97; mem['hE89F]=8'h54;
    mem['hE8A0]=8'h9E; mem['hE8A1]=8'h3B; mem['hE8A2]=8'hBD; mem['hE8A3]=8'hF1;
    mem['hE8A4]=8'h08; mem['hE8A5]=8'hBD; mem['hE8A6]=8'hF3; mem['hE8A7]=8'h79;
    mem['hE8A8]=8'h30; mem['hE8A9]=8'h69; mem['hE8AA]=8'hBD; mem['hE8AB]=8'hF3;
    mem['hE8AC]=8'hDC; mem['hE8AD]=8'hE0; mem['hE8AE]=8'h68; mem['hE8AF]=8'h27;
    mem['hE8B0]=8'h0C; mem['hE8B1]=8'hAE; mem['hE8B2]=8'h6E; mem['hE8B3]=8'h9F;
    mem['hE8B4]=8'h68; mem['hE8B5]=8'hAE; mem['hE8B6]=8'hE8; mem['hE8B7]=8'h10;
    mem['hE8B8]=8'h9F; mem['hE8B9]=8'h83; mem['hE8BA]=8'h7E; mem['hE8BB]=8'hE5;
    mem['hE8BC]=8'h3F; mem['hE8BD]=8'h32; mem['hE8BE]=8'hE8; mem['hE8BF]=8'h12;
    mem['hE8C0]=8'h9D; mem['hE8C1]=8'h82; mem['hE8C2]=8'h81; mem['hE8C3]=8'h2C;
    mem['hE8C4]=8'h26; mem['hE8C5]=8'hF4; mem['hE8C6]=8'h9D; mem['hE8C7]=8'h7C;
    mem['hE8C8]=8'h8D; mem['hE8C9]=8'hBD; mem['hE8CA]=8'h8D; mem['hE8CB]=8'h13;
    mem['hE8CC]=8'h1C; mem['hE8CD]=8'hFE; mem['hE8CE]=8'h7D; mem['hE8CF]=8'h1A;
    mem['hE8D0]=8'h01; mem['hE8D1]=8'h0D; mem['hE8D2]=8'h06; mem['hE8D3]=8'h25;
    mem['hE8D4]=8'h03; mem['hE8D5]=8'h2A; mem['hE8D6]=8'h99; mem['hE8D7]=8'h8C;
    mem['hE8D8]=8'h2B; mem['hE8D9]=8'h96; mem['hE8DA]=8'hC6; mem['hE8DB]=8'h18;
    mem['hE8DC]=8'h7E; mem['hE8DD]=8'hE4; mem['hE8DE]=8'h03; mem['hE8DF]=8'h8D;
    mem['hE8E0]=8'h6E; mem['hE8E1]=8'h4F; mem['hE8E2]=8'h8C; mem['hE8E3]=8'h34;
    mem['hE8E4]=8'h04; mem['hE8E5]=8'h34; mem['hE8E6]=8'h02; mem['hE8E7]=8'hC6;
    mem['hE8E8]=8'h01; mem['hE8E9]=8'hBD; mem['hE8EA]=8'hE3; mem['hE8EB]=8'hF0;
    mem['hE8EC]=8'hBD; mem['hE8ED]=8'hE9; mem['hE8EE]=8'hAC; mem['hE8EF]=8'h0F;
    mem['hE8F0]=8'h3F; mem['hE8F1]=8'h9D; mem['hE8F2]=8'h82; mem['hE8F3]=8'h80;
    mem['hE8F4]=8'hAD; mem['hE8F5]=8'h25; mem['hE8F6]=8'h13; mem['hE8F7]=8'h81;
    mem['hE8F8]=8'h03; mem['hE8F9]=8'h24; mem['hE8FA]=8'h0F; mem['hE8FB]=8'h81;
    mem['hE8FC]=8'h01; mem['hE8FD]=8'h49; mem['hE8FE]=8'h98; mem['hE8FF]=8'h3F;
    mem['hE900]=8'h91; mem['hE901]=8'h3F; mem['hE902]=8'h25; mem['hE903]=8'h64;
    mem['hE904]=8'h97; mem['hE905]=8'h3F; mem['hE906]=8'h9D; mem['hE907]=8'h7C;
    mem['hE908]=8'h20; mem['hE909]=8'hE9; mem['hE90A]=8'hD6; mem['hE90B]=8'h3F;
    mem['hE90C]=8'h26; mem['hE90D]=8'h33; mem['hE90E]=8'h10; mem['hE90F]=8'h24;
    mem['hE910]=8'h00; mem['hE911]=8'h6B; mem['hE912]=8'h8B; mem['hE913]=8'h07;
    mem['hE914]=8'h24; mem['hE915]=8'h67; mem['hE916]=8'h99; mem['hE917]=8'h06;
    mem['hE918]=8'h10; mem['hE919]=8'h27; mem['hE91A]=8'h04; mem['hE91B]=8'h77;
    mem['hE91C]=8'h89; mem['hE91D]=8'hFF; mem['hE91E]=8'h34; mem['hE91F]=8'h02;
    mem['hE920]=8'h48; mem['hE921]=8'hAB; mem['hE922]=8'hE0; mem['hE923]=8'h8E;
    mem['hE924]=8'hE2; mem['hE925]=8'h08; mem['hE926]=8'h30; mem['hE927]=8'h86;
    mem['hE928]=8'h35; mem['hE929]=8'h02; mem['hE92A]=8'hA1; mem['hE92B]=8'h84;
    mem['hE92C]=8'h24; mem['hE92D]=8'h55; mem['hE92E]=8'h8D; mem['hE92F]=8'h9C;
    mem['hE930]=8'h34; mem['hE931]=8'h02; mem['hE932]=8'h8D; mem['hE933]=8'h29;
    mem['hE934]=8'h9E; mem['hE935]=8'h3D; mem['hE936]=8'h35; mem['hE937]=8'h02;
    mem['hE938]=8'h26; mem['hE939]=8'h1D; mem['hE93A]=8'h4D; mem['hE93B]=8'h10;
    mem['hE93C]=8'h27; mem['hE93D]=8'h00; mem['hE93E]=8'h6A; mem['hE93F]=8'h20;
    mem['hE940]=8'h4B; mem['hE941]=8'h08; mem['hE942]=8'h06; mem['hE943]=8'h59;
    mem['hE944]=8'h8D; mem['hE945]=8'h09; mem['hE946]=8'h8E; mem['hE947]=8'hE9;
    mem['hE948]=8'h54; mem['hE949]=8'hD7; mem['hE94A]=8'h3F; mem['hE94B]=8'h0F;
    mem['hE94C]=8'h06; mem['hE94D]=8'h20; mem['hE94E]=8'hD9; mem['hE94F]=8'h9E;
    mem['hE950]=8'h83; mem['hE951]=8'h7E; mem['hE952]=8'hE6; mem['hE953]=8'h68;
    mem['hE954]=8'h64; mem['hE955]=8'hEA; mem['hE956]=8'h78; mem['hE957]=8'hA1;
    mem['hE958]=8'h84; mem['hE959]=8'h24; mem['hE95A]=8'h31; mem['hE95B]=8'h20;
    mem['hE95C]=8'hD3; mem['hE95D]=8'hEC; mem['hE95E]=8'h01; mem['hE95F]=8'h34;
    mem['hE960]=8'h06; mem['hE961]=8'h8D; mem['hE962]=8'h08; mem['hE963]=8'hD6;
    mem['hE964]=8'h3F; mem['hE965]=8'h16; mem['hE966]=8'hFF; mem['hE967]=8'h7B;
    mem['hE968]=8'h7E; mem['hE969]=8'hEA; mem['hE96A]=8'h00; mem['hE96B]=8'hD6;
    mem['hE96C]=8'h54; mem['hE96D]=8'hA6; mem['hE96E]=8'h84; mem['hE96F]=8'h35;
    mem['hE970]=8'h20; mem['hE971]=8'h34; mem['hE972]=8'h04; mem['hE973]=8'hD6;
    mem['hE974]=8'h4F; mem['hE975]=8'h9E; mem['hE976]=8'h50; mem['hE977]=8'hDE;
    mem['hE978]=8'h52; mem['hE979]=8'h34; mem['hE97A]=8'h54; mem['hE97B]=8'h6E;
    mem['hE97C]=8'hA4; mem['hE97D]=8'h9E; mem['hE97E]=8'h74; mem['hE97F]=8'hA6;
    mem['hE980]=8'hE0; mem['hE981]=8'h27; mem['hE982]=8'h26; mem['hE983]=8'h81;
    mem['hE984]=8'h64; mem['hE985]=8'h27; mem['hE986]=8'h03; mem['hE987]=8'hBD;
    mem['hE988]=8'hE8; mem['hE989]=8'hCC; mem['hE98A]=8'h9F; mem['hE98B]=8'h3D;
    mem['hE98C]=8'h35; mem['hE98D]=8'h04; mem['hE98E]=8'h81; mem['hE98F]=8'h5A;
    mem['hE990]=8'h27; mem['hE991]=8'h19; mem['hE992]=8'h81; mem['hE993]=8'h7D;
    mem['hE994]=8'h27; mem['hE995]=8'h15; mem['hE996]=8'h54; mem['hE997]=8'hD7;
    mem['hE998]=8'h0A; mem['hE999]=8'h35; mem['hE99A]=8'h52; mem['hE99B]=8'h97;
    mem['hE99C]=8'h5C; mem['hE99D]=8'h9F; mem['hE99E]=8'h5D; mem['hE99F]=8'hDF;
    mem['hE9A0]=8'h5F; mem['hE9A1]=8'h35; mem['hE9A2]=8'h04; mem['hE9A3]=8'hD7;
    mem['hE9A4]=8'h61; mem['hE9A5]=8'hD8; mem['hE9A6]=8'h54; mem['hE9A7]=8'hD7;
    mem['hE9A8]=8'h62; mem['hE9A9]=8'hD6; mem['hE9AA]=8'h4F; mem['hE9AB]=8'h39;
    mem['hE9AC]=8'hBD; mem['hE9AD]=8'hFB; mem['hE9AE]=8'hF6; mem['hE9AF]=8'h0F;
    mem['hE9B0]=8'h06; mem['hE9B1]=8'h9D; mem['hE9B2]=8'h7C; mem['hE9B3]=8'h24;
    mem['hE9B4]=8'h03; mem['hE9B5]=8'h7E; mem['hE9B6]=8'hF4; mem['hE9B7]=8'h58;
    mem['hE9B8]=8'hBD; mem['hE9B9]=8'hEB; mem['hE9BA]=8'h26; mem['hE9BB]=8'h24;
    mem['hE9BC]=8'h50; mem['hE9BD]=8'h81; mem['hE9BE]=8'h2E; mem['hE9BF]=8'h27;
    mem['hE9C0]=8'hF4; mem['hE9C1]=8'h81; mem['hE9C2]=8'hA7; mem['hE9C3]=8'h27;
    mem['hE9C4]=8'h40; mem['hE9C5]=8'h81; mem['hE9C6]=8'hA6; mem['hE9C7]=8'h27;
    mem['hE9C8]=8'hE3; mem['hE9C9]=8'h81; mem['hE9CA]=8'h22; mem['hE9CB]=8'h26;
    mem['hE9CC]=8'h0A; mem['hE9CD]=8'h9E; mem['hE9CE]=8'h83; mem['hE9CF]=8'hBD;
    mem['hE9D0]=8'hEC; mem['hE9D1]=8'h9C; mem['hE9D2]=8'h9E; mem['hE9D3]=8'h64;
    mem['hE9D4]=8'h9F; mem['hE9D5]=8'h83; mem['hE9D6]=8'h39; mem['hE9D7]=8'h81;
    mem['hE9D8]=8'hA3; mem['hE9D9]=8'h26; mem['hE9DA]=8'h0D; mem['hE9DB]=8'h86;
    mem['hE9DC]=8'h5A; mem['hE9DD]=8'hBD; mem['hE9DE]=8'hE8; mem['hE9DF]=8'hE3;
    mem['hE9E0]=8'hBD; mem['hE9E1]=8'hEB; mem['hE9E2]=8'h71; mem['hE9E3]=8'h43;
    mem['hE9E4]=8'h53; mem['hE9E5]=8'h7E; mem['hE9E6]=8'hEC; mem['hE9E7]=8'h78;
    mem['hE9E8]=8'h4C; mem['hE9E9]=8'h27; mem['hE9EA]=8'h2E; mem['hE9EB]=8'h8D;
    mem['hE9EC]=8'h06; mem['hE9ED]=8'hBD; mem['hE9EE]=8'hE8; mem['hE9EF]=8'hDF;
    mem['hE9F0]=8'hC6; mem['hE9F1]=8'h29; mem['hE9F2]=8'h8C; mem['hE9F3]=8'hC6;
    mem['hE9F4]=8'h28; mem['hE9F5]=8'h8C; mem['hE9F6]=8'hC6; mem['hE9F7]=8'h2C;
    mem['hE9F8]=8'hE1; mem['hE9F9]=8'h9F; mem['hE9FA]=8'h00; mem['hE9FB]=8'h83;
    mem['hE9FC]=8'h26; mem['hE9FD]=8'h02; mem['hE9FE]=8'h0E; mem['hE9FF]=8'h7C;
    mem['hEA00]=8'hC6; mem['hEA01]=8'h02; mem['hEA02]=8'h7E; mem['hEA03]=8'hE4;
    mem['hEA04]=8'h03; mem['hEA05]=8'h86; mem['hEA06]=8'h7D; mem['hEA07]=8'hBD;
    mem['hEA08]=8'hE8; mem['hEA09]=8'hE3; mem['hEA0A]=8'h7E; mem['hEA0B]=8'hF6;
    mem['hEA0C]=8'h2F; mem['hEA0D]=8'hBD; mem['hEA0E]=8'hEA; mem['hEA0F]=8'hDB;
    mem['hEA10]=8'h9F; mem['hEA11]=8'h52; mem['hEA12]=8'h96; mem['hEA13]=8'h06;
    mem['hEA14]=8'h26; mem['hEA15]=8'h95; mem['hEA16]=8'h7E; mem['hEA17]=8'hF3;
    mem['hEA18]=8'h5A; mem['hEA19]=8'h9D; mem['hEA1A]=8'h7C; mem['hEA1B]=8'h1F;
    mem['hEA1C]=8'h89; mem['hEA1D]=8'h58; mem['hEA1E]=8'h9D; mem['hEA1F]=8'h7C;
    mem['hEA20]=8'hC1; mem['hEA21]=8'h38; mem['hEA22]=8'h23; mem['hEA23]=8'h03;
    mem['hEA24]=8'h7E; mem['hEA25]=8'hEA; mem['hEA26]=8'h00; mem['hEA27]=8'h34;
    mem['hEA28]=8'h04; mem['hEA29]=8'hC1; mem['hEA2A]=8'h2A; mem['hEA2B]=8'h25;
    mem['hEA2C]=8'h1E; mem['hEA2D]=8'hC1; mem['hEA2E]=8'h30; mem['hEA2F]=8'h24;
    mem['hEA30]=8'h1C; mem['hEA31]=8'h8D; mem['hEA32]=8'hC0; mem['hEA33]=8'hA6;
    mem['hEA34]=8'hE4; mem['hEA35]=8'hBD; mem['hEA36]=8'hE8; mem['hEA37]=8'hDF;
    mem['hEA38]=8'h8D; mem['hEA39]=8'hBC; mem['hEA3A]=8'hBD; mem['hEA3B]=8'hE8;
    mem['hEA3C]=8'hCF; mem['hEA3D]=8'h35; mem['hEA3E]=8'h02; mem['hEA3F]=8'hDE;
    mem['hEA40]=8'h52; mem['hEA41]=8'h34; mem['hEA42]=8'h42; mem['hEA43]=8'hBD;
    mem['hEA44]=8'hEE; mem['hEA45]=8'h8F; mem['hEA46]=8'h35; mem['hEA47]=8'h02;
    mem['hEA48]=8'h34; mem['hEA49]=8'h06; mem['hEA4A]=8'h8E; mem['hEA4B]=8'h8D;
    mem['hEA4C]=8'h9E; mem['hEA4D]=8'h35; mem['hEA4E]=8'h04; mem['hEA4F]=8'hBE;
    mem['hEA50]=8'hE0; mem['hEA51]=8'hF6; mem['hEA52]=8'h3A; mem['hEA53]=8'hAD;
    mem['hEA54]=8'h94; mem['hEA55]=8'h7E; mem['hEA56]=8'hE8; mem['hEA57]=8'hCC;
    mem['hEA58]=8'h86; mem['hEA59]=8'h4F; mem['hEA5A]=8'h97; mem['hEA5B]=8'h03;
    mem['hEA5C]=8'hBD; mem['hEA5D]=8'hEB; mem['hEA5E]=8'h71; mem['hEA5F]=8'hDD;
    mem['hEA60]=8'h01; mem['hEA61]=8'hBD; mem['hEA62]=8'hF3; mem['hEA63]=8'h90;
    mem['hEA64]=8'hBD; mem['hEA65]=8'hEB; mem['hEA66]=8'h71; mem['hEA67]=8'h0D;
    mem['hEA68]=8'h03; mem['hEA69]=8'h26; mem['hEA6A]=8'h06; mem['hEA6B]=8'h94;
    mem['hEA6C]=8'h01; mem['hEA6D]=8'hD4; mem['hEA6E]=8'h02; mem['hEA6F]=8'h20;
    mem['hEA70]=8'h04; mem['hEA71]=8'h9A; mem['hEA72]=8'h01; mem['hEA73]=8'hDA;
    mem['hEA74]=8'h02; mem['hEA75]=8'h7E; mem['hEA76]=8'hEC; mem['hEA77]=8'h78;
    mem['hEA78]=8'hBD; mem['hEA79]=8'hE8; mem['hEA7A]=8'hD1; mem['hEA7B]=8'h26;
    mem['hEA7C]=8'h10; mem['hEA7D]=8'h96; mem['hEA7E]=8'h61; mem['hEA7F]=8'h8A;
    mem['hEA80]=8'h7F; mem['hEA81]=8'h94; mem['hEA82]=8'h5D; mem['hEA83]=8'h97;
    mem['hEA84]=8'h5D; mem['hEA85]=8'h8E; mem['hEA86]=8'h00; mem['hEA87]=8'h5C;
    mem['hEA88]=8'hBD; mem['hEA89]=8'hF3; mem['hEA8A]=8'hDC; mem['hEA8B]=8'h20;
    mem['hEA8C]=8'h36; mem['hEA8D]=8'h0F; mem['hEA8E]=8'h06; mem['hEA8F]=8'h0A;
    mem['hEA90]=8'h3F; mem['hEA91]=8'hBD; mem['hEA92]=8'hED; mem['hEA93]=8'hDB;
    mem['hEA94]=8'hD7; mem['hEA95]=8'h56; mem['hEA96]=8'h9F; mem['hEA97]=8'h58;
    mem['hEA98]=8'h9E; mem['hEA99]=8'h5F; mem['hEA9A]=8'hBD; mem['hEA9B]=8'hED;
    mem['hEA9C]=8'hDD; mem['hEA9D]=8'h96; mem['hEA9E]=8'h56; mem['hEA9F]=8'h34;
    mem['hEAA0]=8'h04; mem['hEAA1]=8'hA0; mem['hEAA2]=8'hE0; mem['hEAA3]=8'h27;
    mem['hEAA4]=8'h07; mem['hEAA5]=8'h86; mem['hEAA6]=8'h01; mem['hEAA7]=8'h24;
    mem['hEAA8]=8'h03; mem['hEAA9]=8'hD6; mem['hEAAA]=8'h56; mem['hEAAB]=8'h40;
    mem['hEAAC]=8'h97; mem['hEAAD]=8'h54; mem['hEAAE]=8'hDE; mem['hEAAF]=8'h58;
    mem['hEAB0]=8'h5C; mem['hEAB1]=8'h5A; mem['hEAB2]=8'h26; mem['hEAB3]=8'h04;
    mem['hEAB4]=8'hD6; mem['hEAB5]=8'h54; mem['hEAB6]=8'h20; mem['hEAB7]=8'h0B;
    mem['hEAB8]=8'hA6; mem['hEAB9]=8'h80; mem['hEABA]=8'hA1; mem['hEABB]=8'hC0;
    mem['hEABC]=8'h27; mem['hEABD]=8'hF3; mem['hEABE]=8'hC6; mem['hEABF]=8'hFF;
    mem['hEAC0]=8'h24; mem['hEAC1]=8'h01; mem['hEAC2]=8'h50; mem['hEAC3]=8'hCB;
    mem['hEAC4]=8'h01; mem['hEAC5]=8'h59; mem['hEAC6]=8'hD4; mem['hEAC7]=8'h0A;
    mem['hEAC8]=8'h27; mem['hEAC9]=8'h02; mem['hEACA]=8'hC6; mem['hEACB]=8'hFF;
    mem['hEACC]=8'h7E; mem['hEACD]=8'hF3; mem['hEACE]=8'hC2; mem['hEACF]=8'hBD;
    mem['hEAD0]=8'hE9; mem['hEAD1]=8'hF6; mem['hEAD2]=8'hC6; mem['hEAD3]=8'h01;
    mem['hEAD4]=8'h8D; mem['hEAD5]=8'h08; mem['hEAD6]=8'h9D; mem['hEAD7]=8'h82;
    mem['hEAD8]=8'h26; mem['hEAD9]=8'hF5; mem['hEADA]=8'h39; mem['hEADB]=8'h5F;
    mem['hEADC]=8'h9D; mem['hEADD]=8'h82; mem['hEADE]=8'hD7; mem['hEADF]=8'h05;
    mem['hEAE0]=8'h97; mem['hEAE1]=8'h37; mem['hEAE2]=8'h9D; mem['hEAE3]=8'h82;
    mem['hEAE4]=8'h8D; mem['hEAE5]=8'h40; mem['hEAE6]=8'h10; mem['hEAE7]=8'h25;
    mem['hEAE8]=8'hFF; mem['hEAE9]=8'h16; mem['hEAEA]=8'h5F; mem['hEAEB]=8'hD7;
    mem['hEAEC]=8'h06; mem['hEAED]=8'h9D; mem['hEAEE]=8'h7C; mem['hEAEF]=8'h25;
    mem['hEAF0]=8'h04; mem['hEAF1]=8'h8D; mem['hEAF2]=8'h33; mem['hEAF3]=8'h25;
    mem['hEAF4]=8'h0A; mem['hEAF5]=8'h1F; mem['hEAF6]=8'h89; mem['hEAF7]=8'h9D;
    mem['hEAF8]=8'h7C; mem['hEAF9]=8'h25; mem['hEAFA]=8'hFC; mem['hEAFB]=8'h8D;
    mem['hEAFC]=8'h29; mem['hEAFD]=8'h24; mem['hEAFE]=8'hF8; mem['hEAFF]=8'h81;
    mem['hEB00]=8'h24; mem['hEB01]=8'h26; mem['hEB02]=8'h06; mem['hEB03]=8'h03;
    mem['hEB04]=8'h06; mem['hEB05]=8'hCB; mem['hEB06]=8'h80; mem['hEB07]=8'h9D;
    mem['hEB08]=8'h7C; mem['hEB09]=8'hD7; mem['hEB0A]=8'h38; mem['hEB0B]=8'h9A;
    mem['hEB0C]=8'h08; mem['hEB0D]=8'h80; mem['hEB0E]=8'h28; mem['hEB0F]=8'h10;
    mem['hEB10]=8'h27; mem['hEB11]=8'h00; mem['hEB12]=8'h75; mem['hEB13]=8'h0F;
    mem['hEB14]=8'h08; mem['hEB15]=8'h9E; mem['hEB16]=8'h1B; mem['hEB17]=8'hDC;
    mem['hEB18]=8'h37; mem['hEB19]=8'h9C; mem['hEB1A]=8'h1D; mem['hEB1B]=8'h27;
    mem['hEB1C]=8'h12; mem['hEB1D]=8'h10; mem['hEB1E]=8'hA3; mem['hEB1F]=8'h81;
    mem['hEB20]=8'h27; mem['hEB21]=8'h3E; mem['hEB22]=8'h30; mem['hEB23]=8'h05;
    mem['hEB24]=8'h20; mem['hEB25]=8'hF3; mem['hEB26]=8'h81; mem['hEB27]=8'h41;
    mem['hEB28]=8'h25; mem['hEB29]=8'h04; mem['hEB2A]=8'h80; mem['hEB2B]=8'h5B;
    mem['hEB2C]=8'h80; mem['hEB2D]=8'hA5; mem['hEB2E]=8'h39; mem['hEB2F]=8'h8E;
    mem['hEB30]=8'h00; mem['hEB31]=8'h74; mem['hEB32]=8'hEE; mem['hEB33]=8'hE4;
    mem['hEB34]=8'h11; mem['hEB35]=8'h83; mem['hEB36]=8'hEA; mem['hEB37]=8'h10;
    mem['hEB38]=8'h27; mem['hEB39]=8'h28; mem['hEB3A]=8'hDC; mem['hEB3B]=8'h1F;
    mem['hEB3C]=8'hDD; mem['hEB3D]=8'h43; mem['hEB3E]=8'hC3; mem['hEB3F]=8'h00;
    mem['hEB40]=8'h07; mem['hEB41]=8'hDD; mem['hEB42]=8'h41; mem['hEB43]=8'h9E;
    mem['hEB44]=8'h1D; mem['hEB45]=8'h9F; mem['hEB46]=8'h47; mem['hEB47]=8'hBD;
    mem['hEB48]=8'hE3; mem['hEB49]=8'hDB; mem['hEB4A]=8'h9E; mem['hEB4B]=8'h41;
    mem['hEB4C]=8'h9F; mem['hEB4D]=8'h1F; mem['hEB4E]=8'h9E; mem['hEB4F]=8'h45;
    mem['hEB50]=8'h9F; mem['hEB51]=8'h1D; mem['hEB52]=8'h9E; mem['hEB53]=8'h47;
    mem['hEB54]=8'hDC; mem['hEB55]=8'h37; mem['hEB56]=8'hED; mem['hEB57]=8'h81;
    mem['hEB58]=8'h4F; mem['hEB59]=8'h5F; mem['hEB5A]=8'hED; mem['hEB5B]=8'h84;
    mem['hEB5C]=8'hED; mem['hEB5D]=8'h02; mem['hEB5E]=8'hA7; mem['hEB5F]=8'h04;
    mem['hEB60]=8'h9F; mem['hEB61]=8'h39; mem['hEB62]=8'h39; mem['hEB63]=8'h90;
    mem['hEB64]=8'h80; mem['hEB65]=8'h00; mem['hEB66]=8'h00; mem['hEB67]=8'h00;
    mem['hEB68]=8'h9D; mem['hEB69]=8'h7C; mem['hEB6A]=8'hBD; mem['hEB6B]=8'hE8;
    mem['hEB6C]=8'hCA; mem['hEB6D]=8'h96; mem['hEB6E]=8'h54; mem['hEB6F]=8'h2B;
    mem['hEB70]=8'h5D; mem['hEB71]=8'hBD; mem['hEB72]=8'hE8; mem['hEB73]=8'hCC;
    mem['hEB74]=8'h96; mem['hEB75]=8'h4F; mem['hEB76]=8'h81; mem['hEB77]=8'h90;
    mem['hEB78]=8'h25; mem['hEB79]=8'h08; mem['hEB7A]=8'h8E; mem['hEB7B]=8'hEB;
    mem['hEB7C]=8'h63; mem['hEB7D]=8'hBD; mem['hEB7E]=8'hF3; mem['hEB7F]=8'hDC;
    mem['hEB80]=8'h26; mem['hEB81]=8'h4C; mem['hEB82]=8'hBD; mem['hEB83]=8'hF4;
    mem['hEB84]=8'h0E; mem['hEB85]=8'hDC; mem['hEB86]=8'h52; mem['hEB87]=8'h39;
    mem['hEB88]=8'hDC; mem['hEB89]=8'h05; mem['hEB8A]=8'h34; mem['hEB8B]=8'h06;
    mem['hEB8C]=8'h12; mem['hEB8D]=8'h5F; mem['hEB8E]=8'h9E; mem['hEB8F]=8'h37;
    mem['hEB90]=8'h34; mem['hEB91]=8'h14; mem['hEB92]=8'h8D; mem['hEB93]=8'hD4;
    mem['hEB94]=8'h35; mem['hEB95]=8'h34; mem['hEB96]=8'h9F; mem['hEB97]=8'h37;
    mem['hEB98]=8'hDE; mem['hEB99]=8'h52; mem['hEB9A]=8'h34; mem['hEB9B]=8'h60;
    mem['hEB9C]=8'h5C; mem['hEB9D]=8'h9D; mem['hEB9E]=8'h82; mem['hEB9F]=8'h81;
    mem['hEBA0]=8'h2C; mem['hEBA1]=8'h27; mem['hEBA2]=8'hEB; mem['hEBA3]=8'hD7;
    mem['hEBA4]=8'h03; mem['hEBA5]=8'hBD; mem['hEBA6]=8'hE9; mem['hEBA7]=8'hF0;
    mem['hEBA8]=8'h35; mem['hEBA9]=8'h06; mem['hEBAA]=8'hDD; mem['hEBAB]=8'h05;
    mem['hEBAC]=8'h9E; mem['hEBAD]=8'h1D; mem['hEBAE]=8'h9C; mem['hEBAF]=8'h1F;
    mem['hEBB0]=8'h27; mem['hEBB1]=8'h21; mem['hEBB2]=8'hDC; mem['hEBB3]=8'h37;
    mem['hEBB4]=8'h10; mem['hEBB5]=8'hA3; mem['hEBB6]=8'h84; mem['hEBB7]=8'h27;
    mem['hEBB8]=8'h06; mem['hEBB9]=8'hEC; mem['hEBBA]=8'h02; mem['hEBBB]=8'h30;
    mem['hEBBC]=8'h8B; mem['hEBBD]=8'h20; mem['hEBBE]=8'hEF; mem['hEBBF]=8'hC6;
    mem['hEBC0]=8'h12; mem['hEBC1]=8'h96; mem['hEBC2]=8'h05; mem['hEBC3]=8'h26;
    mem['hEBC4]=8'h0B; mem['hEBC5]=8'hD6; mem['hEBC6]=8'h03; mem['hEBC7]=8'hE1;
    mem['hEBC8]=8'h04; mem['hEBC9]=8'h27; mem['hEBCA]=8'h59; mem['hEBCB]=8'hC6;
    mem['hEBCC]=8'h10; mem['hEBCD]=8'h8C; mem['hEBCE]=8'hC6; mem['hEBCF]=8'h08;
    mem['hEBD0]=8'h7E; mem['hEBD1]=8'hE4; mem['hEBD2]=8'h03; mem['hEBD3]=8'hCC;
    mem['hEBD4]=8'h00; mem['hEBD5]=8'h05; mem['hEBD6]=8'hDD; mem['hEBD7]=8'h64;
    mem['hEBD8]=8'hDC; mem['hEBD9]=8'h37; mem['hEBDA]=8'hED; mem['hEBDB]=8'h84;
    mem['hEBDC]=8'hD6; mem['hEBDD]=8'h03; mem['hEBDE]=8'hE7; mem['hEBDF]=8'h04;
    mem['hEBE0]=8'hBD; mem['hEBE1]=8'hE3; mem['hEBE2]=8'hF0; mem['hEBE3]=8'h9F;
    mem['hEBE4]=8'h41; mem['hEBE5]=8'hC6; mem['hEBE6]=8'h0B; mem['hEBE7]=8'h4F;
    mem['hEBE8]=8'h0D; mem['hEBE9]=8'h05; mem['hEBEA]=8'h27; mem['hEBEB]=8'h05;
    mem['hEBEC]=8'h35; mem['hEBED]=8'h06; mem['hEBEE]=8'hC3; mem['hEBEF]=8'h00;
    mem['hEBF0]=8'h01; mem['hEBF1]=8'hED; mem['hEBF2]=8'h05; mem['hEBF3]=8'h8D;
    mem['hEBF4]=8'h5D; mem['hEBF5]=8'hDD; mem['hEBF6]=8'h64; mem['hEBF7]=8'h30;
    mem['hEBF8]=8'h02; mem['hEBF9]=8'h0A; mem['hEBFA]=8'h03; mem['hEBFB]=8'h26;
    mem['hEBFC]=8'hE8; mem['hEBFD]=8'h9F; mem['hEBFE]=8'h0F; mem['hEBFF]=8'hD3;
    mem['hEC00]=8'h0F; mem['hEC01]=8'h10; mem['hEC02]=8'h25; mem['hEC03]=8'hF7;
    mem['hEC04]=8'hFC; mem['hEC05]=8'h1F; mem['hEC06]=8'h01; mem['hEC07]=8'hBD;
    mem['hEC08]=8'hE3; mem['hEC09]=8'hF4; mem['hEC0A]=8'h83; mem['hEC0B]=8'h00;
    mem['hEC0C]=8'h35; mem['hEC0D]=8'hDD; mem['hEC0E]=8'h1F; mem['hEC0F]=8'h4F;
    mem['hEC10]=8'h30; mem['hEC11]=8'h1F; mem['hEC12]=8'hA7; mem['hEC13]=8'h05;
    mem['hEC14]=8'h9C; mem['hEC15]=8'h0F; mem['hEC16]=8'h26; mem['hEC17]=8'hF8;
    mem['hEC18]=8'h9E; mem['hEC19]=8'h41; mem['hEC1A]=8'h96; mem['hEC1B]=8'h1F;
    mem['hEC1C]=8'h93; mem['hEC1D]=8'h41; mem['hEC1E]=8'hED; mem['hEC1F]=8'h02;
    mem['hEC20]=8'h96; mem['hEC21]=8'h05; mem['hEC22]=8'h26; mem['hEC23]=8'h2D;
    mem['hEC24]=8'hE6; mem['hEC25]=8'h04; mem['hEC26]=8'hD7; mem['hEC27]=8'h03;
    mem['hEC28]=8'h4F; mem['hEC29]=8'h5F; mem['hEC2A]=8'hDD; mem['hEC2B]=8'h64;
    mem['hEC2C]=8'h35; mem['hEC2D]=8'h06; mem['hEC2E]=8'hDD; mem['hEC2F]=8'h52;
    mem['hEC30]=8'h10; mem['hEC31]=8'hA3; mem['hEC32]=8'h05; mem['hEC33]=8'h24;
    mem['hEC34]=8'h3A; mem['hEC35]=8'hDE; mem['hEC36]=8'h64; mem['hEC37]=8'h27;
    mem['hEC38]=8'h04; mem['hEC39]=8'h8D; mem['hEC3A]=8'h17; mem['hEC3B]=8'hD3;
    mem['hEC3C]=8'h52; mem['hEC3D]=8'h30; mem['hEC3E]=8'h02; mem['hEC3F]=8'h0A;
    mem['hEC40]=8'h03; mem['hEC41]=8'h26; mem['hEC42]=8'hE7; mem['hEC43]=8'hED;
    mem['hEC44]=8'hE3; mem['hEC45]=8'h58; mem['hEC46]=8'h49; mem['hEC47]=8'h58;
    mem['hEC48]=8'h49; mem['hEC49]=8'hE3; mem['hEC4A]=8'hE1; mem['hEC4B]=8'h30;
    mem['hEC4C]=8'h8B; mem['hEC4D]=8'h30; mem['hEC4E]=8'h05; mem['hEC4F]=8'h9F;
    mem['hEC50]=8'h39; mem['hEC51]=8'h39; mem['hEC52]=8'h86; mem['hEC53]=8'h10;
    mem['hEC54]=8'h97; mem['hEC55]=8'h45; mem['hEC56]=8'hEC; mem['hEC57]=8'h05;
    mem['hEC58]=8'hDD; mem['hEC59]=8'h17; mem['hEC5A]=8'h4F; mem['hEC5B]=8'h5F;
    mem['hEC5C]=8'h58; mem['hEC5D]=8'h49; mem['hEC5E]=8'h25; mem['hEC5F]=8'h0F;
    mem['hEC60]=8'h08; mem['hEC61]=8'h65; mem['hEC62]=8'h09; mem['hEC63]=8'h64;
    mem['hEC64]=8'h24; mem['hEC65]=8'h04; mem['hEC66]=8'hD3; mem['hEC67]=8'h17;
    mem['hEC68]=8'h25; mem['hEC69]=8'h05; mem['hEC6A]=8'h0A; mem['hEC6B]=8'h45;
    mem['hEC6C]=8'h26; mem['hEC6D]=8'hEE; mem['hEC6E]=8'h39; mem['hEC6F]=8'h7E;
    mem['hEC70]=8'hEB; mem['hEC71]=8'hCB; mem['hEC72]=8'h1F; mem['hEC73]=8'h40;
    mem['hEC74]=8'h93; mem['hEC75]=8'h1F; mem['hEC76]=8'h21; mem['hEC77]=8'h4F;
    mem['hEC78]=8'h0F; mem['hEC79]=8'h06; mem['hEC7A]=8'hDD; mem['hEC7B]=8'h50;
    mem['hEC7C]=8'hC6; mem['hEC7D]=8'h90; mem['hEC7E]=8'h7E; mem['hEC7F]=8'hF3;
    mem['hEC80]=8'hC8; mem['hEC81]=8'hBD; mem['hEC82]=8'hE8; mem['hEC83]=8'hCC;
    mem['hEC84]=8'hCE; mem['hEC85]=8'h01; mem['hEC86]=8'hF0; mem['hEC87]=8'hBD;
    mem['hEC88]=8'hF5; mem['hEC89]=8'h22; mem['hEC8A]=8'h32; mem['hEC8B]=8'h62;
    mem['hEC8C]=8'h8E; mem['hEC8D]=8'h01; mem['hEC8E]=8'hEF; mem['hEC8F]=8'h20;
    mem['hEC90]=8'h0B; mem['hEC91]=8'h9F; mem['hEC92]=8'h4D; mem['hEC93]=8'h8D;
    mem['hEC94]=8'h5C; mem['hEC95]=8'h9F; mem['hEC96]=8'h58; mem['hEC97]=8'hD7;
    mem['hEC98]=8'h56; mem['hEC99]=8'h39; mem['hEC9A]=8'h30; mem['hEC9B]=8'h1F;
    mem['hEC9C]=8'h86; mem['hEC9D]=8'h22; mem['hEC9E]=8'h97; mem['hEC9F]=8'h01;
    mem['hECA0]=8'h97; mem['hECA1]=8'h02; mem['hECA2]=8'h30; mem['hECA3]=8'h01;
    mem['hECA4]=8'h9F; mem['hECA5]=8'h62; mem['hECA6]=8'h9F; mem['hECA7]=8'h58;
    mem['hECA8]=8'hC6; mem['hECA9]=8'hFF; mem['hECAA]=8'h5C; mem['hECAB]=8'hA6;
    mem['hECAC]=8'h80; mem['hECAD]=8'h27; mem['hECAE]=8'h0C; mem['hECAF]=8'h91;
    mem['hECB0]=8'h01; mem['hECB1]=8'h27; mem['hECB2]=8'h04; mem['hECB3]=8'h91;
    mem['hECB4]=8'h02; mem['hECB5]=8'h26; mem['hECB6]=8'hF3; mem['hECB7]=8'h81;
    mem['hECB8]=8'h22; mem['hECB9]=8'h27; mem['hECBA]=8'h02; mem['hECBB]=8'h30;
    mem['hECBC]=8'h1F; mem['hECBD]=8'h9F; mem['hECBE]=8'h64; mem['hECBF]=8'hD7;
    mem['hECC0]=8'h56; mem['hECC1]=8'hDE; mem['hECC2]=8'h62; mem['hECC3]=8'h11;
    mem['hECC4]=8'h83; mem['hECC5]=8'h01; mem['hECC6]=8'hF0; mem['hECC7]=8'h22;
    mem['hECC8]=8'h07; mem['hECC9]=8'h8D; mem['hECCA]=8'hC6; mem['hECCB]=8'h9E;
    mem['hECCC]=8'h62; mem['hECCD]=8'hBD; mem['hECCE]=8'hED; mem['hECCF]=8'hC9;
    mem['hECD0]=8'h9E; mem['hECD1]=8'h0B; mem['hECD2]=8'h8C; mem['hECD3]=8'h00;
    mem['hECD4]=8'hF1; mem['hECD5]=8'h26; mem['hECD6]=8'h05; mem['hECD7]=8'hC6;
    mem['hECD8]=8'h1E; mem['hECD9]=8'h7E; mem['hECDA]=8'hE4; mem['hECDB]=8'h03;
    mem['hECDC]=8'h96; mem['hECDD]=8'h56; mem['hECDE]=8'hA7; mem['hECDF]=8'h00;
    mem['hECE0]=8'hDC; mem['hECE1]=8'h58; mem['hECE2]=8'hED; mem['hECE3]=8'h02;
    mem['hECE4]=8'h86; mem['hECE5]=8'hFF; mem['hECE6]=8'h97; mem['hECE7]=8'h06;
    mem['hECE8]=8'h9F; mem['hECE9]=8'h0D; mem['hECEA]=8'h9F; mem['hECEB]=8'h52;
    mem['hECEC]=8'h30; mem['hECED]=8'h05; mem['hECEE]=8'h9F; mem['hECEF]=8'h0B;
    mem['hECF0]=8'h39; mem['hECF1]=8'h0F; mem['hECF2]=8'h07; mem['hECF3]=8'h4F;
    mem['hECF4]=8'h34; mem['hECF5]=8'h06; mem['hECF6]=8'hDC; mem['hECF7]=8'h23;
    mem['hECF8]=8'hA3; mem['hECF9]=8'hE0; mem['hECFA]=8'h10; mem['hECFB]=8'h93;
    mem['hECFC]=8'h21; mem['hECFD]=8'h25; mem['hECFE]=8'h0A; mem['hECFF]=8'hDD;
    mem['hED00]=8'h23; mem['hED01]=8'h9E; mem['hED02]=8'h23; mem['hED03]=8'h30;
    mem['hED04]=8'h01; mem['hED05]=8'h9F; mem['hED06]=8'h25; mem['hED07]=8'h35;
    mem['hED08]=8'h84; mem['hED09]=8'hC6; mem['hED0A]=8'h1A; mem['hED0B]=8'h03;
    mem['hED0C]=8'h07; mem['hED0D]=8'h27; mem['hED0E]=8'hCA; mem['hED0F]=8'h8D;
    mem['hED10]=8'h04; mem['hED11]=8'h35; mem['hED12]=8'h04; mem['hED13]=8'h20;
    mem['hED14]=8'hDE; mem['hED15]=8'h9E; mem['hED16]=8'h27; mem['hED17]=8'h9F;
    mem['hED18]=8'h23; mem['hED19]=8'h4F; mem['hED1A]=8'h5F; mem['hED1B]=8'hDD;
    mem['hED1C]=8'h4B; mem['hED1D]=8'h9E; mem['hED1E]=8'h21; mem['hED1F]=8'h9F;
    mem['hED20]=8'h47; mem['hED21]=8'h8E; mem['hED22]=8'h00; mem['hED23]=8'hC9;
    mem['hED24]=8'h9C; mem['hED25]=8'h0B; mem['hED26]=8'h27; mem['hED27]=8'h04;
    mem['hED28]=8'h8D; mem['hED29]=8'h32; mem['hED2A]=8'h20; mem['hED2B]=8'hF8;
    mem['hED2C]=8'h9E; mem['hED2D]=8'h1B; mem['hED2E]=8'h9C; mem['hED2F]=8'h1D;
    mem['hED30]=8'h27; mem['hED31]=8'h04; mem['hED32]=8'h8D; mem['hED33]=8'h22;
    mem['hED34]=8'h20; mem['hED35]=8'hF8; mem['hED36]=8'h9F; mem['hED37]=8'h41;
    mem['hED38]=8'h9E; mem['hED39]=8'h41; mem['hED3A]=8'h9C; mem['hED3B]=8'h1F;
    mem['hED3C]=8'h27; mem['hED3D]=8'h35; mem['hED3E]=8'hEC; mem['hED3F]=8'h02;
    mem['hED40]=8'hD3; mem['hED41]=8'h41; mem['hED42]=8'hDD; mem['hED43]=8'h41;
    mem['hED44]=8'hA6; mem['hED45]=8'h01; mem['hED46]=8'h2A; mem['hED47]=8'hF0;
    mem['hED48]=8'hE6; mem['hED49]=8'h04; mem['hED4A]=8'h58; mem['hED4B]=8'hCB;
    mem['hED4C]=8'h05; mem['hED4D]=8'h3A; mem['hED4E]=8'h9C; mem['hED4F]=8'h41;
    mem['hED50]=8'h27; mem['hED51]=8'hE8; mem['hED52]=8'h8D; mem['hED53]=8'h08;
    mem['hED54]=8'h20; mem['hED55]=8'hF8; mem['hED56]=8'hA6; mem['hED57]=8'h01;
    mem['hED58]=8'h30; mem['hED59]=8'h02; mem['hED5A]=8'h2A; mem['hED5B]=8'h14;
    mem['hED5C]=8'hE6; mem['hED5D]=8'h84; mem['hED5E]=8'h27; mem['hED5F]=8'h10;
    mem['hED60]=8'hEC; mem['hED61]=8'h02; mem['hED62]=8'h10; mem['hED63]=8'h93;
    mem['hED64]=8'h23; mem['hED65]=8'h22; mem['hED66]=8'h09; mem['hED67]=8'h10;
    mem['hED68]=8'h93; mem['hED69]=8'h47; mem['hED6A]=8'h23; mem['hED6B]=8'h04;
    mem['hED6C]=8'h9F; mem['hED6D]=8'h4B; mem['hED6E]=8'hDD; mem['hED6F]=8'h47;
    mem['hED70]=8'h30; mem['hED71]=8'h05; mem['hED72]=8'h39; mem['hED73]=8'h9E;
    mem['hED74]=8'h4B; mem['hED75]=8'h27; mem['hED76]=8'hFB; mem['hED77]=8'h4F;
    mem['hED78]=8'hE6; mem['hED79]=8'h84; mem['hED7A]=8'h5A; mem['hED7B]=8'hD3;
    mem['hED7C]=8'h47; mem['hED7D]=8'hDD; mem['hED7E]=8'h43; mem['hED7F]=8'h9E;
    mem['hED80]=8'h23; mem['hED81]=8'h9F; mem['hED82]=8'h41; mem['hED83]=8'hBD;
    mem['hED84]=8'hE3; mem['hED85]=8'hDD; mem['hED86]=8'h9E; mem['hED87]=8'h4B;
    mem['hED88]=8'hDC; mem['hED89]=8'h45; mem['hED8A]=8'hED; mem['hED8B]=8'h02;
    mem['hED8C]=8'h9E; mem['hED8D]=8'h45; mem['hED8E]=8'h30; mem['hED8F]=8'h1F;
    mem['hED90]=8'h7E; mem['hED91]=8'hED; mem['hED92]=8'h17; mem['hED93]=8'hDC;
    mem['hED94]=8'h52; mem['hED95]=8'h34; mem['hED96]=8'h06; mem['hED97]=8'hBD;
    mem['hED98]=8'hE9; mem['hED99]=8'hAC; mem['hED9A]=8'hBD; mem['hED9B]=8'hE8;
    mem['hED9C]=8'hCF; mem['hED9D]=8'h35; mem['hED9E]=8'h10; mem['hED9F]=8'h9F;
    mem['hEDA0]=8'h62; mem['hEDA1]=8'hE6; mem['hEDA2]=8'h84; mem['hEDA3]=8'h9E;
    mem['hEDA4]=8'h52; mem['hEDA5]=8'hEB; mem['hEDA6]=8'h84; mem['hEDA7]=8'h24;
    mem['hEDA8]=8'h05; mem['hEDA9]=8'hC6; mem['hEDAA]=8'h1C; mem['hEDAB]=8'h7E;
    mem['hEDAC]=8'hE4; mem['hEDAD]=8'h03; mem['hEDAE]=8'hBD; mem['hEDAF]=8'hEC;
    mem['hEDB0]=8'h91; mem['hEDB1]=8'h9E; mem['hEDB2]=8'h62; mem['hEDB3]=8'hE6;
    mem['hEDB4]=8'h84; mem['hEDB5]=8'h8D; mem['hEDB6]=8'h10; mem['hEDB7]=8'h9E;
    mem['hEDB8]=8'h4D; mem['hEDB9]=8'h8D; mem['hEDBA]=8'h22; mem['hEDBB]=8'h8D;
    mem['hEDBC]=8'h0C; mem['hEDBD]=8'h9E; mem['hEDBE]=8'h62; mem['hEDBF]=8'h8D;
    mem['hEDC0]=8'h1C; mem['hEDC1]=8'hBD; mem['hEDC2]=8'hEC; mem['hEDC3]=8'hD0;
    mem['hEDC4]=8'h7E; mem['hEDC5]=8'hE8; mem['hEDC6]=8'hF1; mem['hEDC7]=8'hAE;
    mem['hEDC8]=8'h02; mem['hEDC9]=8'hDE; mem['hEDCA]=8'h25; mem['hEDCB]=8'h5C;
    mem['hEDCC]=8'h20; mem['hEDCD]=8'h04; mem['hEDCE]=8'hA6; mem['hEDCF]=8'h80;
    mem['hEDD0]=8'hA7; mem['hEDD1]=8'hC0; mem['hEDD2]=8'h5A; mem['hEDD3]=8'h26;
    mem['hEDD4]=8'hF9; mem['hEDD5]=8'hDF; mem['hEDD6]=8'h25; mem['hEDD7]=8'h39;
    mem['hEDD8]=8'hBD; mem['hEDD9]=8'hE8; mem['hEDDA]=8'hCF; mem['hEDDB]=8'h9E;
    mem['hEDDC]=8'h52; mem['hEDDD]=8'hE6; mem['hEDDE]=8'h84; mem['hEDDF]=8'h8D;
    mem['hEDE0]=8'h18; mem['hEDE1]=8'h26; mem['hEDE2]=8'h13; mem['hEDE3]=8'hAE;
    mem['hEDE4]=8'h07; mem['hEDE5]=8'h30; mem['hEDE6]=8'h1F; mem['hEDE7]=8'h9C;
    mem['hEDE8]=8'h23; mem['hEDE9]=8'h26; mem['hEDEA]=8'h08; mem['hEDEB]=8'h34;
    mem['hEDEC]=8'h04; mem['hEDED]=8'hD3; mem['hEDEE]=8'h23; mem['hEDEF]=8'hDD;
    mem['hEDF0]=8'h23; mem['hEDF1]=8'h35; mem['hEDF2]=8'h04; mem['hEDF3]=8'h30;
    mem['hEDF4]=8'h01; mem['hEDF5]=8'h39; mem['hEDF6]=8'hAE; mem['hEDF7]=8'h02;
    mem['hEDF8]=8'h39; mem['hEDF9]=8'h9C; mem['hEDFA]=8'h0D; mem['hEDFB]=8'h26;
    mem['hEDFC]=8'h07; mem['hEDFD]=8'h9F; mem['hEDFE]=8'h0B; mem['hEDFF]=8'h30;
    mem['hEE00]=8'h1B; mem['hEE01]=8'h9F; mem['hEE02]=8'h0D; mem['hEE03]=8'h4F;
    mem['hEE04]=8'h39; mem['hEE05]=8'h8D; mem['hEE06]=8'h03; mem['hEE07]=8'h7E;
    mem['hEE08]=8'hEC; mem['hEE09]=8'h77; mem['hEE0A]=8'h8D; mem['hEE0B]=8'hCC;
    mem['hEE0C]=8'h0F; mem['hEE0D]=8'h06; mem['hEE0E]=8'h5D; mem['hEE0F]=8'h39;
    mem['hEE10]=8'hBD; mem['hEE11]=8'hEE; mem['hEE12]=8'h92; mem['hEE13]=8'hC6;
    mem['hEE14]=8'h01; mem['hEE15]=8'hBD; mem['hEE16]=8'hEC; mem['hEE17]=8'hF1;
    mem['hEE18]=8'h96; mem['hEE19]=8'h53; mem['hEE1A]=8'hBD; mem['hEE1B]=8'hEC;
    mem['hEE1C]=8'h95; mem['hEE1D]=8'hA7; mem['hEE1E]=8'h84; mem['hEE1F]=8'h32;
    mem['hEE20]=8'h62; mem['hEE21]=8'h7E; mem['hEE22]=8'hEC; mem['hEE23]=8'hD0;
    mem['hEE24]=8'h8D; mem['hEE25]=8'h02; mem['hEE26]=8'h20; mem['hEE27]=8'hDF;
    mem['hEE28]=8'h8D; mem['hEE29]=8'hE0; mem['hEE2A]=8'h27; mem['hEE2B]=8'h5E;
    mem['hEE2C]=8'hE6; mem['hEE2D]=8'h84; mem['hEE2E]=8'h39; mem['hEE2F]=8'h8D;
    mem['hEE30]=8'h48; mem['hEE31]=8'h4F; mem['hEE32]=8'hE1; mem['hEE33]=8'h84;
    mem['hEE34]=8'h23; mem['hEE35]=8'h03; mem['hEE36]=8'hE6; mem['hEE37]=8'h84;
    mem['hEE38]=8'h4F; mem['hEE39]=8'h34; mem['hEE3A]=8'h06; mem['hEE3B]=8'hBD;
    mem['hEE3C]=8'hEC; mem['hEE3D]=8'h93; mem['hEE3E]=8'h9E; mem['hEE3F]=8'h4D;
    mem['hEE40]=8'h8D; mem['hEE41]=8'h9B; mem['hEE42]=8'h35; mem['hEE43]=8'h04;
    mem['hEE44]=8'h3A; mem['hEE45]=8'h35; mem['hEE46]=8'h04; mem['hEE47]=8'hBD;
    mem['hEE48]=8'hED; mem['hEE49]=8'hC9; mem['hEE4A]=8'h20; mem['hEE4B]=8'hD5;
    mem['hEE4C]=8'h8D; mem['hEE4D]=8'h2B; mem['hEE4E]=8'hA0; mem['hEE4F]=8'h84;
    mem['hEE50]=8'h40; mem['hEE51]=8'h20; mem['hEE52]=8'hDF; mem['hEE53]=8'hC6;
    mem['hEE54]=8'hFF; mem['hEE55]=8'hD7; mem['hEE56]=8'h53; mem['hEE57]=8'h9D;
    mem['hEE58]=8'h82; mem['hEE59]=8'h81; mem['hEE5A]=8'h29; mem['hEE5B]=8'h27;
    mem['hEE5C]=8'h05; mem['hEE5D]=8'hBD; mem['hEE5E]=8'hE9; mem['hEE5F]=8'hF6;
    mem['hEE60]=8'h8D; mem['hEE61]=8'h2D; mem['hEE62]=8'h8D; mem['hEE63]=8'h15;
    mem['hEE64]=8'h27; mem['hEE65]=8'h24; mem['hEE66]=8'h5F; mem['hEE67]=8'h4A;
    mem['hEE68]=8'hA1; mem['hEE69]=8'h84; mem['hEE6A]=8'h24; mem['hEE6B]=8'hCD;
    mem['hEE6C]=8'h1F; mem['hEE6D]=8'h89; mem['hEE6E]=8'hE0; mem['hEE6F]=8'h84;
    mem['hEE70]=8'h50; mem['hEE71]=8'hD1; mem['hEE72]=8'h53; mem['hEE73]=8'h23;
    mem['hEE74]=8'hC4; mem['hEE75]=8'hD6; mem['hEE76]=8'h53; mem['hEE77]=8'h20;
    mem['hEE78]=8'hC0; mem['hEE79]=8'hBD; mem['hEE7A]=8'hE9; mem['hEE7B]=8'hF0;
    mem['hEE7C]=8'hEE; mem['hEE7D]=8'hE4; mem['hEE7E]=8'hAE; mem['hEE7F]=8'h65;
    mem['hEE80]=8'h9F; mem['hEE81]=8'h4D; mem['hEE82]=8'hA6; mem['hEE83]=8'h64;
    mem['hEE84]=8'hE6; mem['hEE85]=8'h64; mem['hEE86]=8'h32; mem['hEE87]=8'h67;
    mem['hEE88]=8'h1F; mem['hEE89]=8'h35; mem['hEE8A]=8'h7E; mem['hEE8B]=8'hEB;
    mem['hEE8C]=8'hCE; mem['hEE8D]=8'h9D; mem['hEE8E]=8'h7C; mem['hEE8F]=8'hBD;
    mem['hEE90]=8'hE8; mem['hEE91]=8'hCA; mem['hEE92]=8'hBD; mem['hEE93]=8'hEB;
    mem['hEE94]=8'h6D; mem['hEE95]=8'h4D; mem['hEE96]=8'h26; mem['hEE97]=8'hF2;
    mem['hEE98]=8'h0E; mem['hEE99]=8'h82; mem['hEE9A]=8'hBD; mem['hEE9B]=8'hEE;
    mem['hEE9C]=8'h0A; mem['hEE9D]=8'h10; mem['hEE9E]=8'h27; mem['hEE9F]=8'h02;
    mem['hEEA0]=8'hDE; mem['hEEA1]=8'hDE; mem['hEEA2]=8'h83; mem['hEEA3]=8'h9F;
    mem['hEEA4]=8'h83; mem['hEEA5]=8'h3A; mem['hEEA6]=8'hA6; mem['hEEA7]=8'h84;
    mem['hEEA8]=8'h34; mem['hEEA9]=8'h52; mem['hEEAA]=8'h6F; mem['hEEAB]=8'h84;
    mem['hEEAC]=8'h9D; mem['hEEAD]=8'h82; mem['hEEAE]=8'hBD; mem['hEEAF]=8'hF4;
    mem['hEEB0]=8'h58; mem['hEEB1]=8'h35; mem['hEEB2]=8'h52; mem['hEEB3]=8'hA7;
    mem['hEEB4]=8'h84; mem['hEEB5]=8'hDF; mem['hEEB6]=8'h83; mem['hEEB7]=8'h39;
    mem['hEEB8]=8'h8D; mem['hEEB9]=8'h07; mem['hEEBA]=8'h9F; mem['hEEBB]=8'h2B;
    mem['hEEBC]=8'hBD; mem['hEEBD]=8'hE9; mem['hEEBE]=8'hF6; mem['hEEBF]=8'h20;
    mem['hEEC0]=8'hCE; mem['hEEC1]=8'hBD; mem['hEEC2]=8'hE8; mem['hEEC3]=8'hCA;
    mem['hEEC4]=8'h96; mem['hEEC5]=8'h54; mem['hEEC6]=8'h2B; mem['hEEC7]=8'hC2;
    mem['hEEC8]=8'h96; mem['hEEC9]=8'h4F; mem['hEECA]=8'h81; mem['hEECB]=8'h90;
    mem['hEECC]=8'h22; mem['hEECD]=8'hBC; mem['hEECE]=8'hBD; mem['hEECF]=8'hF4;
    mem['hEED0]=8'h0E; mem['hEED1]=8'h9E; mem['hEED2]=8'h52; mem['hEED3]=8'h39;
    mem['hEED4]=8'h8D; mem['hEED5]=8'hEE; mem['hEED6]=8'hE6; mem['hEED7]=8'h84;
    mem['hEED8]=8'h7E; mem['hEED9]=8'hEC; mem['hEEDA]=8'h77; mem['hEEDB]=8'h8D;
    mem['hEEDC]=8'hDB; mem['hEEDD]=8'h9E; mem['hEEDE]=8'h2B; mem['hEEDF]=8'hE7;
    mem['hEEE0]=8'h84; mem['hEEE1]=8'h39; mem['hEEE2]=8'h34; mem['hEEE3]=8'h01;
    mem['hEEE4]=8'hBD; mem['hEEE5]=8'hE7; mem['hEEE6]=8'h14; mem['hEEE7]=8'hBD;
    mem['hEEE8]=8'hE4; mem['hEEE9]=8'hA2; mem['hEEEA]=8'h9F; mem['hEEEB]=8'h66;
    mem['hEEEC]=8'h35; mem['hEEED]=8'h01; mem['hEEEE]=8'h27; mem['hEEEF]=8'h12;
    mem['hEEF0]=8'h9D; mem['hEEF1]=8'h82; mem['hEEF2]=8'h27; mem['hEEF3]=8'h13;
    mem['hEEF4]=8'h81; mem['hEEF5]=8'hA7; mem['hEEF6]=8'h26; mem['hEEF7]=8'h09;
    mem['hEEF8]=8'h9D; mem['hEEF9]=8'h7C; mem['hEEFA]=8'h27; mem['hEEFB]=8'h06;
    mem['hEEFC]=8'hBD; mem['hEEFD]=8'hE7; mem['hEEFE]=8'h14; mem['hEEFF]=8'h27;
    mem['hEF00]=8'h06; mem['hEF01]=8'h39; mem['hEF02]=8'hCE; mem['hEF03]=8'hFF;
    mem['hEF04]=8'hFF; mem['hEF05]=8'hDF; mem['hEF06]=8'h2B; mem['hEF07]=8'h32;
    mem['hEF08]=8'h62; mem['hEF09]=8'h9E; mem['hEF0A]=8'h66; mem['hEF0B]=8'hBD;
    mem['hEF0C]=8'hF0; mem['hEF0D]=8'hA6; mem['hEF0E]=8'hBD; mem['hEF0F]=8'hE1;
    mem['hEF10]=8'h97; mem['hEF11]=8'hEC; mem['hEF12]=8'h84; mem['hEF13]=8'h26;
    mem['hEF14]=8'h03; mem['hEF15]=8'h7E; mem['hEF16]=8'hE4; mem['hEF17]=8'h22;
    mem['hEF18]=8'h9F; mem['hEF19]=8'h66; mem['hEF1A]=8'hEC; mem['hEF1B]=8'h02;
    mem['hEF1C]=8'h10; mem['hEF1D]=8'h93; mem['hEF1E]=8'h2B; mem['hEF1F]=8'h22;
    mem['hEF20]=8'hF4; mem['hEF21]=8'hBD; mem['hEF22]=8'hF5; mem['hEF23]=8'h12;
    mem['hEF24]=8'hBD; mem['hEF25]=8'hF0; mem['hEF26]=8'hF2; mem['hEF27]=8'h9E;
    mem['hEF28]=8'h66; mem['hEF29]=8'h8D; mem['hEF2A]=8'h10; mem['hEF2B]=8'hAE;
    mem['hEF2C]=8'h9F; mem['hEF2D]=8'h00; mem['hEF2E]=8'h66; mem['hEF2F]=8'hCE;
    mem['hEF30]=8'h00; mem['hEF31]=8'hF4; mem['hEF32]=8'hA6; mem['hEF33]=8'hC0;
    mem['hEF34]=8'h27; mem['hEF35]=8'hD5; mem['hEF36]=8'hBD; mem['hEF37]=8'hF0;
    mem['hEF38]=8'hF7; mem['hEF39]=8'h20; mem['hEF3A]=8'hF7; mem['hEF3B]=8'h30;
    mem['hEF3C]=8'h04; mem['hEF3D]=8'h10; mem['hEF3E]=8'h8E; mem['hEF3F]=8'h00;
    mem['hEF40]=8'hF4; mem['hEF41]=8'hA6; mem['hEF42]=8'h80; mem['hEF43]=8'h27;
    mem['hEF44]=8'h51; mem['hEF45]=8'h2B; mem['hEF46]=8'h15; mem['hEF47]=8'h81;
    mem['hEF48]=8'h3A; mem['hEF49]=8'h26; mem['hEF4A]=8'h0D; mem['hEF4B]=8'hE6;
    mem['hEF4C]=8'h84; mem['hEF4D]=8'hC1; mem['hEF4E]=8'h84; mem['hEF4F]=8'h27;
    mem['hEF50]=8'hF0; mem['hEF51]=8'hC1; mem['hEF52]=8'h83; mem['hEF53]=8'h27;
    mem['hEF54]=8'hEC; mem['hEF55]=8'h8C; mem['hEF56]=8'h86; mem['hEF57]=8'h21;
    mem['hEF58]=8'h8D; mem['hEF59]=8'h30; mem['hEF5A]=8'h20; mem['hEF5B]=8'hE5;
    mem['hEF5C]=8'hCE; mem['hEF5D]=8'hE0; mem['hEF5E]=8'hE4; mem['hEF5F]=8'h81;
    mem['hEF60]=8'hFF; mem['hEF61]=8'h26; mem['hEF62]=8'h04; mem['hEF63]=8'hA6;
    mem['hEF64]=8'h80; mem['hEF65]=8'h33; mem['hEF66]=8'h45; mem['hEF67]=8'h84;
    mem['hEF68]=8'h7F; mem['hEF69]=8'h33; mem['hEF6A]=8'h4A; mem['hEF6B]=8'h6D;
    mem['hEF6C]=8'hC4; mem['hEF6D]=8'h27; mem['hEF6E]=8'hE7; mem['hEF6F]=8'hA0;
    mem['hEF70]=8'hC4; mem['hEF71]=8'h2A; mem['hEF72]=8'hF6; mem['hEF73]=8'hAB;
    mem['hEF74]=8'hC4; mem['hEF75]=8'hEE; mem['hEF76]=8'h41; mem['hEF77]=8'h4A;
    mem['hEF78]=8'h2B; mem['hEF79]=8'h06; mem['hEF7A]=8'h6D; mem['hEF7B]=8'hC0;
    mem['hEF7C]=8'h2A; mem['hEF7D]=8'hFC; mem['hEF7E]=8'h20; mem['hEF7F]=8'hF7;
    mem['hEF80]=8'hA6; mem['hEF81]=8'hC4; mem['hEF82]=8'h8D; mem['hEF83]=8'h06;
    mem['hEF84]=8'h6D; mem['hEF85]=8'hC0; mem['hEF86]=8'h2A; mem['hEF87]=8'hF8;
    mem['hEF88]=8'h20; mem['hEF89]=8'hB7; mem['hEF8A]=8'h10; mem['hEF8B]=8'h8C;
    mem['hEF8C]=8'h01; mem['hEF8D]=8'hED; mem['hEF8E]=8'h24; mem['hEF8F]=8'h06;
    mem['hEF90]=8'h84; mem['hEF91]=8'h7F; mem['hEF92]=8'hA7; mem['hEF93]=8'hA0;
    mem['hEF94]=8'h6F; mem['hEF95]=8'hA4; mem['hEF96]=8'h39; mem['hEF97]=8'h9E;
    mem['hEF98]=8'h83; mem['hEF99]=8'hCE; mem['hEF9A]=8'h00; mem['hEF9B]=8'hF3;
    mem['hEF9C]=8'h0F; mem['hEF9D]=8'h43; mem['hEF9E]=8'h0F; mem['hEF9F]=8'h44;
    mem['hEFA0]=8'hA6; mem['hEFA1]=8'h80; mem['hEFA2]=8'h27; mem['hEFA3]=8'h21;
    mem['hEFA4]=8'h0D; mem['hEFA5]=8'h43; mem['hEFA6]=8'h27; mem['hEFA7]=8'h0F;
    mem['hEFA8]=8'hBD; mem['hEFA9]=8'hEB; mem['hEFAA]=8'h26; mem['hEFAB]=8'h24;
    mem['hEFAC]=8'h18; mem['hEFAD]=8'h81; mem['hEFAE]=8'h30; mem['hEFAF]=8'h25;
    mem['hEFB0]=8'h04; mem['hEFB1]=8'h81; mem['hEFB2]=8'h39; mem['hEFB3]=8'h23;
    mem['hEFB4]=8'h10; mem['hEFB5]=8'h0F; mem['hEFB6]=8'h43; mem['hEFB7]=8'h81;
    mem['hEFB8]=8'h20; mem['hEFB9]=8'h27; mem['hEFBA]=8'h0A; mem['hEFBB]=8'h97;
    mem['hEFBC]=8'h42; mem['hEFBD]=8'h81; mem['hEFBE]=8'h22; mem['hEFBF]=8'h27;
    mem['hEFC0]=8'h38; mem['hEFC1]=8'h0D; mem['hEFC2]=8'h44; mem['hEFC3]=8'h27;
    mem['hEFC4]=8'h19; mem['hEFC5]=8'hA7; mem['hEFC6]=8'hC0; mem['hEFC7]=8'h27;
    mem['hEFC8]=8'h06; mem['hEFC9]=8'h81; mem['hEFCA]=8'h3A; mem['hEFCB]=8'h27;
    mem['hEFCC]=8'hCF; mem['hEFCD]=8'h20; mem['hEFCE]=8'hD1; mem['hEFCF]=8'h6F;
    mem['hEFD0]=8'hC0; mem['hEFD1]=8'h6F; mem['hEFD2]=8'hC0; mem['hEFD3]=8'h1F;
    mem['hEFD4]=8'h30; mem['hEFD5]=8'h83; mem['hEFD6]=8'h00; mem['hEFD7]=8'hF1;
    mem['hEFD8]=8'h8E; mem['hEFD9]=8'h00; mem['hEFDA]=8'hF2; mem['hEFDB]=8'h9F;
    mem['hEFDC]=8'h83; mem['hEFDD]=8'h39; mem['hEFDE]=8'h81; mem['hEFDF]=8'h3F;
    mem['hEFE0]=8'h26; mem['hEFE1]=8'h04; mem['hEFE2]=8'h86; mem['hEFE3]=8'h87;
    mem['hEFE4]=8'h20; mem['hEFE5]=8'hDF; mem['hEFE6]=8'h81; mem['hEFE7]=8'h27;
    mem['hEFE8]=8'h26; mem['hEFE9]=8'h13; mem['hEFEA]=8'hCC; mem['hEFEB]=8'h3A;
    mem['hEFEC]=8'h83; mem['hEFED]=8'hED; mem['hEFEE]=8'hC1; mem['hEFEF]=8'h0F;
    mem['hEFF0]=8'h42; mem['hEFF1]=8'hA6; mem['hEFF2]=8'h80; mem['hEFF3]=8'h27;
    mem['hEFF4]=8'hD0; mem['hEFF5]=8'h91; mem['hEFF6]=8'h42; mem['hEFF7]=8'h27;
    mem['hEFF8]=8'hCC; mem['hEFF9]=8'hA7; mem['hEFFA]=8'hC0; mem['hEFFB]=8'h20;
    mem['hEFFC]=8'hF4; mem['hEFFD]=8'h81; mem['hEFFE]=8'h30; mem['hEFFF]=8'h25;
    mem['hF000]=8'h04; mem['hF001]=8'h81; mem['hF002]=8'h3C; mem['hF003]=8'h25;
    mem['hF004]=8'hC0; mem['hF005]=8'h30; mem['hF006]=8'h1F; mem['hF007]=8'h34;
    mem['hF008]=8'h50; mem['hF009]=8'h0F; mem['hF00A]=8'h41; mem['hF00B]=8'hCE;
    mem['hF00C]=8'hE0; mem['hF00D]=8'hE4; mem['hF00E]=8'h0F; mem['hF00F]=8'h42;
    mem['hF010]=8'h33; mem['hF011]=8'h4A; mem['hF012]=8'hA6; mem['hF013]=8'hC4;
    mem['hF014]=8'h27; mem['hF015]=8'h31; mem['hF016]=8'h10; mem['hF017]=8'hAE;
    mem['hF018]=8'h41; mem['hF019]=8'hAE; mem['hF01A]=8'hE4; mem['hF01B]=8'hE6;
    mem['hF01C]=8'hA0; mem['hF01D]=8'hE0; mem['hF01E]=8'h80; mem['hF01F]=8'h27;
    mem['hF020]=8'hFA; mem['hF021]=8'hC1; mem['hF022]=8'h80; mem['hF023]=8'h26;
    mem['hF024]=8'h38; mem['hF025]=8'h32; mem['hF026]=8'h62; mem['hF027]=8'h35;
    mem['hF028]=8'h40; mem['hF029]=8'hDA; mem['hF02A]=8'h42; mem['hF02B]=8'h96;
    mem['hF02C]=8'h41; mem['hF02D]=8'h26; mem['hF02E]=8'h06; mem['hF02F]=8'hC1;
    mem['hF030]=8'h84; mem['hF031]=8'h26; mem['hF032]=8'h06; mem['hF033]=8'h86;
    mem['hF034]=8'h3A; mem['hF035]=8'hED; mem['hF036]=8'hC1; mem['hF037]=8'h20;
    mem['hF038]=8'h94; mem['hF039]=8'hE7; mem['hF03A]=8'hC0; mem['hF03B]=8'hC1;
    mem['hF03C]=8'h86; mem['hF03D]=8'h26; mem['hF03E]=8'h02; mem['hF03F]=8'h0C;
    mem['hF040]=8'h44; mem['hF041]=8'hC1; mem['hF042]=8'h82; mem['hF043]=8'h27;
    mem['hF044]=8'hAA; mem['hF045]=8'h20; mem['hF046]=8'h86; mem['hF047]=8'hCE;
    mem['hF048]=8'hE0; mem['hF049]=8'hE9; mem['hF04A]=8'h03; mem['hF04B]=8'h41;
    mem['hF04C]=8'h26; mem['hF04D]=8'hC0; mem['hF04E]=8'h35; mem['hF04F]=8'h50;
    mem['hF050]=8'hA6; mem['hF051]=8'h80; mem['hF052]=8'hA7; mem['hF053]=8'hC0;
    mem['hF054]=8'hBD; mem['hF055]=8'hEB; mem['hF056]=8'h26; mem['hF057]=8'h25;
    mem['hF058]=8'hEC; mem['hF059]=8'h03; mem['hF05A]=8'h43; mem['hF05B]=8'h20;
    mem['hF05C]=8'hE8; mem['hF05D]=8'h0C; mem['hF05E]=8'h42; mem['hF05F]=8'h4A;
    mem['hF060]=8'h27; mem['hF061]=8'hAE; mem['hF062]=8'h31; mem['hF063]=8'h3F;
    mem['hF064]=8'hE6; mem['hF065]=8'hA0; mem['hF066]=8'h2A; mem['hF067]=8'hFC;
    mem['hF068]=8'h20; mem['hF069]=8'hAF; mem['hF06A]=8'h27; mem['hF06B]=8'h36;
    mem['hF06C]=8'h8D; mem['hF06D]=8'h01; mem['hF06E]=8'h39; mem['hF06F]=8'h27;
    mem['hF070]=8'h3E; mem['hF071]=8'h81; mem['hF072]=8'h9F; mem['hF073]=8'h27;
    mem['hF074]=8'h53; mem['hF075]=8'h81; mem['hF076]=8'h2C; mem['hF077]=8'h27;
    mem['hF078]=8'h37; mem['hF079]=8'h81; mem['hF07A]=8'h3B; mem['hF07B]=8'h27;
    mem['hF07C]=8'h60; mem['hF07D]=8'hBD; mem['hF07E]=8'hE8; mem['hF07F]=8'hDF;
    mem['hF080]=8'h96; mem['hF081]=8'h06; mem['hF082]=8'h34; mem['hF083]=8'h02;
    mem['hF084]=8'h26; mem['hF085]=8'h06; mem['hF086]=8'hBD; mem['hF087]=8'hF5;
    mem['hF088]=8'h1F; mem['hF089]=8'hBD; mem['hF08A]=8'hEC; mem['hF08B]=8'h9A;
    mem['hF08C]=8'h8D; mem['hF08D]=8'h57; mem['hF08E]=8'h35; mem['hF08F]=8'h04;
    mem['hF090]=8'hBD; mem['hF091]=8'hE1; mem['hF092]=8'h30; mem['hF093]=8'h5D;
    mem['hF094]=8'h26; mem['hF095]=8'h08; mem['hF096]=8'h9D; mem['hF097]=8'h82;
    mem['hF098]=8'h81; mem['hF099]=8'h2C; mem['hF09A]=8'h27; mem['hF09B]=8'h14;
    mem['hF09C]=8'h8D; mem['hF09D]=8'h54; mem['hF09E]=8'h9D; mem['hF09F]=8'h82;
    mem['hF0A0]=8'h26; mem['hF0A1]=8'hCF; mem['hF0A2]=8'h86; mem['hF0A3]=8'h0D;
    mem['hF0A4]=8'h20; mem['hF0A5]=8'h51; mem['hF0A6]=8'hBD; mem['hF0A7]=8'hE1;
    mem['hF0A8]=8'h30; mem['hF0A9]=8'h27; mem['hF0AA]=8'hF7; mem['hF0AB]=8'h96;
    mem['hF0AC]=8'h6C; mem['hF0AD]=8'h26; mem['hF0AE]=8'hF3; mem['hF0AF]=8'h39;
    mem['hF0B0]=8'hBD; mem['hF0B1]=8'hE1; mem['hF0B2]=8'h30; mem['hF0B3]=8'h27;
    mem['hF0B4]=8'h0A; mem['hF0B5]=8'hD6; mem['hF0B6]=8'h6C; mem['hF0B7]=8'hD1;
    mem['hF0B8]=8'h6B; mem['hF0B9]=8'h25; mem['hF0BA]=8'h06; mem['hF0BB]=8'h8D;
    mem['hF0BC]=8'hE5; mem['hF0BD]=8'h20; mem['hF0BE]=8'h1E; mem['hF0BF]=8'hD6;
    mem['hF0C0]=8'h6C; mem['hF0C1]=8'hD0; mem['hF0C2]=8'h6A; mem['hF0C3]=8'h24;
    mem['hF0C4]=8'hFC; mem['hF0C5]=8'h50; mem['hF0C6]=8'h20; mem['hF0C7]=8'h10;
    mem['hF0C8]=8'hBD; mem['hF0C9]=8'hEE; mem['hF0CA]=8'h8D; mem['hF0CB]=8'h81;
    mem['hF0CC]=8'h29; mem['hF0CD]=8'h10; mem['hF0CE]=8'h26; mem['hF0CF]=8'hF9;
    mem['hF0D0]=8'h2F; mem['hF0D1]=8'hBD; mem['hF0D2]=8'hE1; mem['hF0D3]=8'h30;
    mem['hF0D4]=8'hD0; mem['hF0D5]=8'h6C; mem['hF0D6]=8'h23; mem['hF0D7]=8'h05;
    mem['hF0D8]=8'h8D; mem['hF0D9]=8'h18; mem['hF0DA]=8'h5A; mem['hF0DB]=8'h26;
    mem['hF0DC]=8'hFB; mem['hF0DD]=8'h9D; mem['hF0DE]=8'h7C; mem['hF0DF]=8'h7E;
    mem['hF0E0]=8'hF0; mem['hF0E1]=8'h6F; mem['hF0E2]=8'hBD; mem['hF0E3]=8'hEC;
    mem['hF0E4]=8'h9C; mem['hF0E5]=8'hBD; mem['hF0E6]=8'hED; mem['hF0E7]=8'hDB;
    mem['hF0E8]=8'h5C; mem['hF0E9]=8'h5A; mem['hF0EA]=8'h27; mem['hF0EB]=8'hC3;
    mem['hF0EC]=8'hA6; mem['hF0ED]=8'h80; mem['hF0EE]=8'h8D; mem['hF0EF]=8'h07;
    mem['hF0F0]=8'h20; mem['hF0F1]=8'hF7; mem['hF0F2]=8'h86; mem['hF0F3]=8'h20;
    mem['hF0F4]=8'h8C; mem['hF0F5]=8'h86; mem['hF0F6]=8'h3F; mem['hF0F7]=8'h7E;
    mem['hF0F8]=8'hE0; mem['hF0F9]=8'h14; mem['hF0FA]=8'h8E; mem['hF0FB]=8'hF6;
    mem['hF0FC]=8'h06; mem['hF0FD]=8'h20; mem['hF0FE]=8'h09; mem['hF0FF]=8'hBD;
    mem['hF100]=8'hF2; mem['hF101]=8'h75; mem['hF102]=8'h03; mem['hF103]=8'h54;
    mem['hF104]=8'h03; mem['hF105]=8'h62; mem['hF106]=8'h20; mem['hF107]=8'h03;
    mem['hF108]=8'hBD; mem['hF109]=8'hF2; mem['hF10A]=8'h75; mem['hF10B]=8'h5D;
    mem['hF10C]=8'h10; mem['hF10D]=8'h27; mem['hF10E]=8'h02; mem['hF10F]=8'h80;
    mem['hF110]=8'h8E; mem['hF111]=8'h00; mem['hF112]=8'h5C; mem['hF113]=8'h1F;
    mem['hF114]=8'h89; mem['hF115]=8'h5D; mem['hF116]=8'h27; mem['hF117]=8'h6C;
    mem['hF118]=8'hD0; mem['hF119]=8'h4F; mem['hF11A]=8'h27; mem['hF11B]=8'h69;
    mem['hF11C]=8'h25; mem['hF11D]=8'h0A; mem['hF11E]=8'h97; mem['hF11F]=8'h4F;
    mem['hF120]=8'h96; mem['hF121]=8'h61; mem['hF122]=8'h97; mem['hF123]=8'h54;
    mem['hF124]=8'h8E; mem['hF125]=8'h00; mem['hF126]=8'h4F; mem['hF127]=8'h50;
    mem['hF128]=8'hC1; mem['hF129]=8'hF8; mem['hF12A]=8'h2F; mem['hF12B]=8'h59;
    mem['hF12C]=8'h4F; mem['hF12D]=8'h64; mem['hF12E]=8'h01; mem['hF12F]=8'hBD;
    mem['hF130]=8'hF2; mem['hF131]=8'h00; mem['hF132]=8'hD6; mem['hF133]=8'h62;
    mem['hF134]=8'h2A; mem['hF135]=8'h0B; mem['hF136]=8'h63; mem['hF137]=8'h01;
    mem['hF138]=8'h63; mem['hF139]=8'h02; mem['hF13A]=8'h63; mem['hF13B]=8'h03;
    mem['hF13C]=8'h63; mem['hF13D]=8'h04; mem['hF13E]=8'h43; mem['hF13F]=8'h89;
    mem['hF140]=8'h00; mem['hF141]=8'h97; mem['hF142]=8'h63; mem['hF143]=8'h96;
    mem['hF144]=8'h53; mem['hF145]=8'h99; mem['hF146]=8'h60; mem['hF147]=8'h97;
    mem['hF148]=8'h53; mem['hF149]=8'h96; mem['hF14A]=8'h52; mem['hF14B]=8'h99;
    mem['hF14C]=8'h5F; mem['hF14D]=8'h97; mem['hF14E]=8'h52; mem['hF14F]=8'h96;
    mem['hF150]=8'h51; mem['hF151]=8'h99; mem['hF152]=8'h5E; mem['hF153]=8'h97;
    mem['hF154]=8'h51; mem['hF155]=8'h96; mem['hF156]=8'h50; mem['hF157]=8'h99;
    mem['hF158]=8'h5D; mem['hF159]=8'h97; mem['hF15A]=8'h50; mem['hF15B]=8'h5D;
    mem['hF15C]=8'h2A; mem['hF15D]=8'h44; mem['hF15E]=8'h25; mem['hF15F]=8'h02;
    mem['hF160]=8'h8D; mem['hF161]=8'h5D; mem['hF162]=8'h5F; mem['hF163]=8'h96;
    mem['hF164]=8'h50; mem['hF165]=8'h26; mem['hF166]=8'h2E; mem['hF167]=8'h96;
    mem['hF168]=8'h51; mem['hF169]=8'h97; mem['hF16A]=8'h50; mem['hF16B]=8'h96;
    mem['hF16C]=8'h52; mem['hF16D]=8'h97; mem['hF16E]=8'h51; mem['hF16F]=8'h96;
    mem['hF170]=8'h53; mem['hF171]=8'h97; mem['hF172]=8'h52; mem['hF173]=8'h96;
    mem['hF174]=8'h63; mem['hF175]=8'h97; mem['hF176]=8'h53; mem['hF177]=8'h0F;
    mem['hF178]=8'h63; mem['hF179]=8'hCB; mem['hF17A]=8'h08; mem['hF17B]=8'hC1;
    mem['hF17C]=8'h28; mem['hF17D]=8'h2D; mem['hF17E]=8'hE4; mem['hF17F]=8'h4F;
    mem['hF180]=8'h97; mem['hF181]=8'h4F; mem['hF182]=8'h97; mem['hF183]=8'h54;
    mem['hF184]=8'h39; mem['hF185]=8'h8D; mem['hF186]=8'h6D; mem['hF187]=8'h5F;
    mem['hF188]=8'h20; mem['hF189]=8'hA8; mem['hF18A]=8'h5C; mem['hF18B]=8'h08;
    mem['hF18C]=8'h63; mem['hF18D]=8'h09; mem['hF18E]=8'h53; mem['hF18F]=8'h09;
    mem['hF190]=8'h52; mem['hF191]=8'h09; mem['hF192]=8'h51; mem['hF193]=8'h09;
    mem['hF194]=8'h50; mem['hF195]=8'h2A; mem['hF196]=8'hF3; mem['hF197]=8'h96;
    mem['hF198]=8'h4F; mem['hF199]=8'h34; mem['hF19A]=8'h04; mem['hF19B]=8'hA0;
    mem['hF19C]=8'hE0; mem['hF19D]=8'h97; mem['hF19E]=8'h4F; mem['hF19F]=8'h23;
    mem['hF1A0]=8'hDE; mem['hF1A1]=8'h8C; mem['hF1A2]=8'h25; mem['hF1A3]=8'h08;
    mem['hF1A4]=8'h08; mem['hF1A5]=8'h63; mem['hF1A6]=8'h86; mem['hF1A7]=8'h00;
    mem['hF1A8]=8'h97; mem['hF1A9]=8'h63; mem['hF1AA]=8'h20; mem['hF1AB]=8'h0C;
    mem['hF1AC]=8'h0C; mem['hF1AD]=8'h4F; mem['hF1AE]=8'h27; mem['hF1AF]=8'h28;
    mem['hF1B0]=8'h06; mem['hF1B1]=8'h50; mem['hF1B2]=8'h06; mem['hF1B3]=8'h51;
    mem['hF1B4]=8'h06; mem['hF1B5]=8'h52; mem['hF1B6]=8'h06; mem['hF1B7]=8'h53;
    mem['hF1B8]=8'h24; mem['hF1B9]=8'h04; mem['hF1BA]=8'h8D; mem['hF1BB]=8'h0D;
    mem['hF1BC]=8'h27; mem['hF1BD]=8'hEE; mem['hF1BE]=8'h39; mem['hF1BF]=8'h03;
    mem['hF1C0]=8'h54; mem['hF1C1]=8'h03; mem['hF1C2]=8'h50; mem['hF1C3]=8'h03;
    mem['hF1C4]=8'h51; mem['hF1C5]=8'h03; mem['hF1C6]=8'h52; mem['hF1C7]=8'h03;
    mem['hF1C8]=8'h53; mem['hF1C9]=8'h9E; mem['hF1CA]=8'h52; mem['hF1CB]=8'h30;
    mem['hF1CC]=8'h01; mem['hF1CD]=8'h9F; mem['hF1CE]=8'h52; mem['hF1CF]=8'h26;
    mem['hF1D0]=8'h06; mem['hF1D1]=8'h9E; mem['hF1D2]=8'h50; mem['hF1D3]=8'h30;
    mem['hF1D4]=8'h01; mem['hF1D5]=8'h9F; mem['hF1D6]=8'h50; mem['hF1D7]=8'h39;
    mem['hF1D8]=8'hC6; mem['hF1D9]=8'h0A; mem['hF1DA]=8'h7E; mem['hF1DB]=8'hE4;
    mem['hF1DC]=8'h03; mem['hF1DD]=8'h8E; mem['hF1DE]=8'h00; mem['hF1DF]=8'h12;
    mem['hF1E0]=8'hA6; mem['hF1E1]=8'h04; mem['hF1E2]=8'h97; mem['hF1E3]=8'h63;
    mem['hF1E4]=8'hA6; mem['hF1E5]=8'h03; mem['hF1E6]=8'hA7; mem['hF1E7]=8'h04;
    mem['hF1E8]=8'hA6; mem['hF1E9]=8'h02; mem['hF1EA]=8'hA7; mem['hF1EB]=8'h03;
    mem['hF1EC]=8'hA6; mem['hF1ED]=8'h01; mem['hF1EE]=8'hA7; mem['hF1EF]=8'h02;
    mem['hF1F0]=8'h96; mem['hF1F1]=8'h5B; mem['hF1F2]=8'hA7; mem['hF1F3]=8'h01;
    mem['hF1F4]=8'hCB; mem['hF1F5]=8'h08; mem['hF1F6]=8'h2F; mem['hF1F7]=8'hE8;
    mem['hF1F8]=8'h96; mem['hF1F9]=8'h63; mem['hF1FA]=8'hC0; mem['hF1FB]=8'h08;
    mem['hF1FC]=8'h27; mem['hF1FD]=8'h0C; mem['hF1FE]=8'h67; mem['hF1FF]=8'h01;
    mem['hF200]=8'h66; mem['hF201]=8'h02; mem['hF202]=8'h66; mem['hF203]=8'h03;
    mem['hF204]=8'h66; mem['hF205]=8'h04; mem['hF206]=8'h46; mem['hF207]=8'h5C;
    mem['hF208]=8'h26; mem['hF209]=8'hF4; mem['hF20A]=8'h39; mem['hF20B]=8'h81;
    mem['hF20C]=8'h00; mem['hF20D]=8'h00; mem['hF20E]=8'h00; mem['hF20F]=8'h00;
    mem['hF210]=8'h8D; mem['hF211]=8'h63; mem['hF212]=8'h27; mem['hF213]=8'h60;
    mem['hF214]=8'h8D; mem['hF215]=8'h78; mem['hF216]=8'h86; mem['hF217]=8'h00;
    mem['hF218]=8'h97; mem['hF219]=8'h13; mem['hF21A]=8'h97; mem['hF21B]=8'h14;
    mem['hF21C]=8'h97; mem['hF21D]=8'h15; mem['hF21E]=8'h97; mem['hF21F]=8'h16;
    mem['hF220]=8'hD6; mem['hF221]=8'h53; mem['hF222]=8'h8D; mem['hF223]=8'h22;
    mem['hF224]=8'hD6; mem['hF225]=8'h63; mem['hF226]=8'hD7; mem['hF227]=8'h8B;
    mem['hF228]=8'hD6; mem['hF229]=8'h52; mem['hF22A]=8'h8D; mem['hF22B]=8'h1A;
    mem['hF22C]=8'hD6; mem['hF22D]=8'h63; mem['hF22E]=8'hD7; mem['hF22F]=8'h8A;
    mem['hF230]=8'hD6; mem['hF231]=8'h51; mem['hF232]=8'h8D; mem['hF233]=8'h12;
    mem['hF234]=8'hD6; mem['hF235]=8'h63; mem['hF236]=8'hD7; mem['hF237]=8'h89;
    mem['hF238]=8'hD6; mem['hF239]=8'h50; mem['hF23A]=8'h8D; mem['hF23B]=8'h0C;
    mem['hF23C]=8'hD6; mem['hF23D]=8'h63; mem['hF23E]=8'hD7; mem['hF23F]=8'h88;
    mem['hF240]=8'hBD; mem['hF241]=8'hF3; mem['hF242]=8'h51; mem['hF243]=8'h7E;
    mem['hF244]=8'hF1; mem['hF245]=8'h62; mem['hF246]=8'h27; mem['hF247]=8'h95;
    mem['hF248]=8'h43; mem['hF249]=8'h96; mem['hF24A]=8'h13; mem['hF24B]=8'h56;
    mem['hF24C]=8'h27; mem['hF24D]=8'h26; mem['hF24E]=8'h24; mem['hF24F]=8'h16;
    mem['hF250]=8'h96; mem['hF251]=8'h16; mem['hF252]=8'h9B; mem['hF253]=8'h60;
    mem['hF254]=8'h97; mem['hF255]=8'h16; mem['hF256]=8'h96; mem['hF257]=8'h15;
    mem['hF258]=8'h99; mem['hF259]=8'h5F; mem['hF25A]=8'h97; mem['hF25B]=8'h15;
    mem['hF25C]=8'h96; mem['hF25D]=8'h14; mem['hF25E]=8'h99; mem['hF25F]=8'h5E;
    mem['hF260]=8'h97; mem['hF261]=8'h14; mem['hF262]=8'h96; mem['hF263]=8'h13;
    mem['hF264]=8'h99; mem['hF265]=8'h5D; mem['hF266]=8'h46; mem['hF267]=8'h97;
    mem['hF268]=8'h13; mem['hF269]=8'h06; mem['hF26A]=8'h14; mem['hF26B]=8'h06;
    mem['hF26C]=8'h15; mem['hF26D]=8'h06; mem['hF26E]=8'h16; mem['hF26F]=8'h06;
    mem['hF270]=8'h63; mem['hF271]=8'h4F; mem['hF272]=8'h20; mem['hF273]=8'hD5;
    mem['hF274]=8'h39; mem['hF275]=8'hEC; mem['hF276]=8'h01; mem['hF277]=8'h97;
    mem['hF278]=8'h61; mem['hF279]=8'h8A; mem['hF27A]=8'h80; mem['hF27B]=8'hDD;
    mem['hF27C]=8'h5D; mem['hF27D]=8'hD6; mem['hF27E]=8'h61; mem['hF27F]=8'hD8;
    mem['hF280]=8'h54; mem['hF281]=8'hD7; mem['hF282]=8'h62; mem['hF283]=8'hEC;
    mem['hF284]=8'h03; mem['hF285]=8'hDD; mem['hF286]=8'h5F; mem['hF287]=8'hA6;
    mem['hF288]=8'h84; mem['hF289]=8'h97; mem['hF28A]=8'h5C; mem['hF28B]=8'hD6;
    mem['hF28C]=8'h4F; mem['hF28D]=8'h39; mem['hF28E]=8'h4D; mem['hF28F]=8'h27;
    mem['hF290]=8'h16; mem['hF291]=8'h9B; mem['hF292]=8'h4F; mem['hF293]=8'h46;
    mem['hF294]=8'h49; mem['hF295]=8'h28; mem['hF296]=8'h10; mem['hF297]=8'h8B;
    mem['hF298]=8'h80; mem['hF299]=8'h97; mem['hF29A]=8'h4F; mem['hF29B]=8'h27;
    mem['hF29C]=8'h0C; mem['hF29D]=8'h96; mem['hF29E]=8'h62; mem['hF29F]=8'h97;
    mem['hF2A0]=8'h54; mem['hF2A1]=8'h39; mem['hF2A2]=8'h96; mem['hF2A3]=8'h54;
    mem['hF2A4]=8'h43; mem['hF2A5]=8'h20; mem['hF2A6]=8'h02; mem['hF2A7]=8'h32;
    mem['hF2A8]=8'h62; mem['hF2A9]=8'h10; mem['hF2AA]=8'h2A; mem['hF2AB]=8'hFE;
    mem['hF2AC]=8'hD2; mem['hF2AD]=8'h7E; mem['hF2AE]=8'hF1; mem['hF2AF]=8'hD8;
    mem['hF2B0]=8'hBD; mem['hF2B1]=8'hF3; mem['hF2B2]=8'hA5; mem['hF2B3]=8'h27;
    mem['hF2B4]=8'h0D; mem['hF2B5]=8'h8B; mem['hF2B6]=8'h02; mem['hF2B7]=8'h25;
    mem['hF2B8]=8'hF4; mem['hF2B9]=8'h0F; mem['hF2BA]=8'h62; mem['hF2BB]=8'hBD;
    mem['hF2BC]=8'hF1; mem['hF2BD]=8'h13; mem['hF2BE]=8'h0C; mem['hF2BF]=8'h4F;
    mem['hF2C0]=8'h27; mem['hF2C1]=8'hEB; mem['hF2C2]=8'h39; mem['hF2C3]=8'h84;
    mem['hF2C4]=8'h20; mem['hF2C5]=8'h00; mem['hF2C6]=8'h00; mem['hF2C7]=8'h00;
    mem['hF2C8]=8'hBD; mem['hF2C9]=8'hF3; mem['hF2CA]=8'hA5; mem['hF2CB]=8'h8E;
    mem['hF2CC]=8'hF2; mem['hF2CD]=8'hC3; mem['hF2CE]=8'h5F; mem['hF2CF]=8'hD7;
    mem['hF2D0]=8'h62; mem['hF2D1]=8'hBD; mem['hF2D2]=8'hF3; mem['hF2D3]=8'h5A;
    mem['hF2D4]=8'h8C; mem['hF2D5]=8'h8D; mem['hF2D6]=8'h9E; mem['hF2D7]=8'h27;
    mem['hF2D8]=8'h73; mem['hF2D9]=8'h00; mem['hF2DA]=8'h4F; mem['hF2DB]=8'h8D;
    mem['hF2DC]=8'hB1; mem['hF2DD]=8'h0C; mem['hF2DE]=8'h4F; mem['hF2DF]=8'h27;
    mem['hF2E0]=8'hCC; mem['hF2E1]=8'h8E; mem['hF2E2]=8'h00; mem['hF2E3]=8'h13;
    mem['hF2E4]=8'hC6; mem['hF2E5]=8'h04; mem['hF2E6]=8'hD7; mem['hF2E7]=8'h03;
    mem['hF2E8]=8'hC6; mem['hF2E9]=8'h01; mem['hF2EA]=8'h96; mem['hF2EB]=8'h50;
    mem['hF2EC]=8'h91; mem['hF2ED]=8'h5D; mem['hF2EE]=8'h26; mem['hF2EF]=8'h13;
    mem['hF2F0]=8'h96; mem['hF2F1]=8'h51; mem['hF2F2]=8'h91; mem['hF2F3]=8'h5E;
    mem['hF2F4]=8'h26; mem['hF2F5]=8'h0D; mem['hF2F6]=8'h96; mem['hF2F7]=8'h52;
    mem['hF2F8]=8'h91; mem['hF2F9]=8'h5F; mem['hF2FA]=8'h26; mem['hF2FB]=8'h07;
    mem['hF2FC]=8'h96; mem['hF2FD]=8'h53; mem['hF2FE]=8'h91; mem['hF2FF]=8'h60;
    mem['hF300]=8'h26; mem['hF301]=8'h01; mem['hF302]=8'h43; mem['hF303]=8'h1F;
    mem['hF304]=8'hA8; mem['hF305]=8'h59; mem['hF306]=8'h24; mem['hF307]=8'h0A;
    mem['hF308]=8'hE7; mem['hF309]=8'h80; mem['hF30A]=8'h0A; mem['hF30B]=8'h03;
    mem['hF30C]=8'h2B; mem['hF30D]=8'h34; mem['hF30E]=8'h27; mem['hF30F]=8'h2E;
    mem['hF310]=8'hC6; mem['hF311]=8'h01; mem['hF312]=8'h1F; mem['hF313]=8'h8A;
    mem['hF314]=8'h25; mem['hF315]=8'h0E; mem['hF316]=8'h08; mem['hF317]=8'h60;
    mem['hF318]=8'h09; mem['hF319]=8'h5F; mem['hF31A]=8'h09; mem['hF31B]=8'h5E;
    mem['hF31C]=8'h09; mem['hF31D]=8'h5D; mem['hF31E]=8'h25; mem['hF31F]=8'hE3;
    mem['hF320]=8'h2B; mem['hF321]=8'hC8; mem['hF322]=8'h20; mem['hF323]=8'hDF;
    mem['hF324]=8'h96; mem['hF325]=8'h60; mem['hF326]=8'h90; mem['hF327]=8'h53;
    mem['hF328]=8'h97; mem['hF329]=8'h60; mem['hF32A]=8'h96; mem['hF32B]=8'h5F;
    mem['hF32C]=8'h92; mem['hF32D]=8'h52; mem['hF32E]=8'h97; mem['hF32F]=8'h5F;
    mem['hF330]=8'h96; mem['hF331]=8'h5E; mem['hF332]=8'h92; mem['hF333]=8'h51;
    mem['hF334]=8'h97; mem['hF335]=8'h5E; mem['hF336]=8'h96; mem['hF337]=8'h5D;
    mem['hF338]=8'h92; mem['hF339]=8'h50; mem['hF33A]=8'h97; mem['hF33B]=8'h5D;
    mem['hF33C]=8'h20; mem['hF33D]=8'hD8; mem['hF33E]=8'hC6; mem['hF33F]=8'h40;
    mem['hF340]=8'h20; mem['hF341]=8'hD0; mem['hF342]=8'h56; mem['hF343]=8'h56;
    mem['hF344]=8'h56; mem['hF345]=8'hD7; mem['hF346]=8'h63; mem['hF347]=8'h8D;
    mem['hF348]=8'h08; mem['hF349]=8'h7E; mem['hF34A]=8'hF1; mem['hF34B]=8'h62;
    mem['hF34C]=8'hC6; mem['hF34D]=8'h14; mem['hF34E]=8'h7E; mem['hF34F]=8'hE4;
    mem['hF350]=8'h03; mem['hF351]=8'h9E; mem['hF352]=8'h13; mem['hF353]=8'h9F;
    mem['hF354]=8'h50; mem['hF355]=8'h9E; mem['hF356]=8'h15; mem['hF357]=8'h9F;
    mem['hF358]=8'h52; mem['hF359]=8'h39; mem['hF35A]=8'h34; mem['hF35B]=8'h02;
    mem['hF35C]=8'hEC; mem['hF35D]=8'h01; mem['hF35E]=8'h97; mem['hF35F]=8'h54;
    mem['hF360]=8'h8A; mem['hF361]=8'h80; mem['hF362]=8'hDD; mem['hF363]=8'h50;
    mem['hF364]=8'h0F; mem['hF365]=8'h63; mem['hF366]=8'hE6; mem['hF367]=8'h84;
    mem['hF368]=8'hAE; mem['hF369]=8'h03; mem['hF36A]=8'h9F; mem['hF36B]=8'h52;
    mem['hF36C]=8'hD7; mem['hF36D]=8'h4F; mem['hF36E]=8'h35; mem['hF36F]=8'h82;
    mem['hF370]=8'h8E; mem['hF371]=8'h00; mem['hF372]=8'h45; mem['hF373]=8'h20;
    mem['hF374]=8'h06; mem['hF375]=8'h8E; mem['hF376]=8'h00; mem['hF377]=8'h40;
    mem['hF378]=8'h8C; mem['hF379]=8'h9E; mem['hF37A]=8'h3B; mem['hF37B]=8'h96;
    mem['hF37C]=8'h4F; mem['hF37D]=8'hA7; mem['hF37E]=8'h84; mem['hF37F]=8'h96;
    mem['hF380]=8'h54; mem['hF381]=8'h8A; mem['hF382]=8'h7F; mem['hF383]=8'h94;
    mem['hF384]=8'h50; mem['hF385]=8'hA7; mem['hF386]=8'h01; mem['hF387]=8'h96;
    mem['hF388]=8'h51; mem['hF389]=8'hA7; mem['hF38A]=8'h02; mem['hF38B]=8'hDE;
    mem['hF38C]=8'h52; mem['hF38D]=8'hEF; mem['hF38E]=8'h03; mem['hF38F]=8'h39;
    mem['hF390]=8'h96; mem['hF391]=8'h61; mem['hF392]=8'h97; mem['hF393]=8'h54;
    mem['hF394]=8'h9E; mem['hF395]=8'h5C; mem['hF396]=8'h9F; mem['hF397]=8'h4F;
    mem['hF398]=8'h0F; mem['hF399]=8'h63; mem['hF39A]=8'h96; mem['hF39B]=8'h5E;
    mem['hF39C]=8'h97; mem['hF39D]=8'h51; mem['hF39E]=8'h96; mem['hF39F]=8'h54;
    mem['hF3A0]=8'h9E; mem['hF3A1]=8'h5F; mem['hF3A2]=8'h9F; mem['hF3A3]=8'h52;
    mem['hF3A4]=8'h39; mem['hF3A5]=8'hDC; mem['hF3A6]=8'h4F; mem['hF3A7]=8'hDD;
    mem['hF3A8]=8'h5C; mem['hF3A9]=8'h9E; mem['hF3AA]=8'h51; mem['hF3AB]=8'h9F;
    mem['hF3AC]=8'h5E; mem['hF3AD]=8'h9E; mem['hF3AE]=8'h53; mem['hF3AF]=8'h9F;
    mem['hF3B0]=8'h60; mem['hF3B1]=8'h4D; mem['hF3B2]=8'h39; mem['hF3B3]=8'hD6;
    mem['hF3B4]=8'h4F; mem['hF3B5]=8'h27; mem['hF3B6]=8'h08; mem['hF3B7]=8'hD6;
    mem['hF3B8]=8'h54; mem['hF3B9]=8'h59; mem['hF3BA]=8'hC6; mem['hF3BB]=8'hFF;
    mem['hF3BC]=8'h25; mem['hF3BD]=8'h01; mem['hF3BE]=8'h50; mem['hF3BF]=8'h39;
    mem['hF3C0]=8'h8D; mem['hF3C1]=8'hF1; mem['hF3C2]=8'hD7; mem['hF3C3]=8'h50;
    mem['hF3C4]=8'h0F; mem['hF3C5]=8'h51; mem['hF3C6]=8'hC6; mem['hF3C7]=8'h88;
    mem['hF3C8]=8'h96; mem['hF3C9]=8'h50; mem['hF3CA]=8'h80; mem['hF3CB]=8'h80;
    mem['hF3CC]=8'hD7; mem['hF3CD]=8'h4F; mem['hF3CE]=8'hDC; mem['hF3CF]=8'h74;
    mem['hF3D0]=8'hDD; mem['hF3D1]=8'h52; mem['hF3D2]=8'h97; mem['hF3D3]=8'h63;
    mem['hF3D4]=8'h97; mem['hF3D5]=8'h54; mem['hF3D6]=8'h7E; mem['hF3D7]=8'hF1;
    mem['hF3D8]=8'h5E; mem['hF3D9]=8'h0F; mem['hF3DA]=8'h54; mem['hF3DB]=8'h39;
    mem['hF3DC]=8'hE6; mem['hF3DD]=8'h84; mem['hF3DE]=8'h27; mem['hF3DF]=8'hD3;
    mem['hF3E0]=8'hE6; mem['hF3E1]=8'h01; mem['hF3E2]=8'hD8; mem['hF3E3]=8'h54;
    mem['hF3E4]=8'h2B; mem['hF3E5]=8'hD1; mem['hF3E6]=8'hD6; mem['hF3E7]=8'h4F;
    mem['hF3E8]=8'hE1; mem['hF3E9]=8'h84; mem['hF3EA]=8'h26; mem['hF3EB]=8'h1D;
    mem['hF3EC]=8'hE6; mem['hF3ED]=8'h01; mem['hF3EE]=8'hCA; mem['hF3EF]=8'h7F;
    mem['hF3F0]=8'hD4; mem['hF3F1]=8'h50; mem['hF3F2]=8'hE1; mem['hF3F3]=8'h01;
    mem['hF3F4]=8'h26; mem['hF3F5]=8'h13; mem['hF3F6]=8'hD6; mem['hF3F7]=8'h51;
    mem['hF3F8]=8'hE1; mem['hF3F9]=8'h02; mem['hF3FA]=8'h26; mem['hF3FB]=8'h0D;
    mem['hF3FC]=8'hD6; mem['hF3FD]=8'h52; mem['hF3FE]=8'hE1; mem['hF3FF]=8'h03;
    mem['hF400]=8'h26; mem['hF401]=8'h07; mem['hF402]=8'hD6; mem['hF403]=8'h53;
    mem['hF404]=8'hE0; mem['hF405]=8'h04; mem['hF406]=8'h26; mem['hF407]=8'h01;
    mem['hF408]=8'h39; mem['hF409]=8'h56; mem['hF40A]=8'hD8; mem['hF40B]=8'h54;
    mem['hF40C]=8'h20; mem['hF40D]=8'hAB; mem['hF40E]=8'hD6; mem['hF40F]=8'h4F;
    mem['hF410]=8'h27; mem['hF411]=8'h3D; mem['hF412]=8'hC0; mem['hF413]=8'hA0;
    mem['hF414]=8'h96; mem['hF415]=8'h54; mem['hF416]=8'h2A; mem['hF417]=8'h05;
    mem['hF418]=8'h03; mem['hF419]=8'h5B; mem['hF41A]=8'hBD; mem['hF41B]=8'hF1;
    mem['hF41C]=8'hC1; mem['hF41D]=8'h8E; mem['hF41E]=8'h00; mem['hF41F]=8'h4F;
    mem['hF420]=8'hC1; mem['hF421]=8'hF8; mem['hF422]=8'h2E; mem['hF423]=8'h06;
    mem['hF424]=8'hBD; mem['hF425]=8'hF1; mem['hF426]=8'hF4; mem['hF427]=8'h0F;
    mem['hF428]=8'h5B; mem['hF429]=8'h39; mem['hF42A]=8'h0F; mem['hF42B]=8'h5B;
    mem['hF42C]=8'h96; mem['hF42D]=8'h54; mem['hF42E]=8'h49; mem['hF42F]=8'h06;
    mem['hF430]=8'h50; mem['hF431]=8'h7E; mem['hF432]=8'hF2; mem['hF433]=8'h00;
    mem['hF434]=8'hD6; mem['hF435]=8'h4F; mem['hF436]=8'hC1; mem['hF437]=8'hA0;
    mem['hF438]=8'h24; mem['hF439]=8'h1D; mem['hF43A]=8'h8D; mem['hF43B]=8'hD2;
    mem['hF43C]=8'hD7; mem['hF43D]=8'h63; mem['hF43E]=8'h96; mem['hF43F]=8'h54;
    mem['hF440]=8'hD7; mem['hF441]=8'h54; mem['hF442]=8'h80; mem['hF443]=8'h80;
    mem['hF444]=8'h86; mem['hF445]=8'hA0; mem['hF446]=8'h97; mem['hF447]=8'h4F;
    mem['hF448]=8'h96; mem['hF449]=8'h53; mem['hF44A]=8'h97; mem['hF44B]=8'h01;
    mem['hF44C]=8'h7E; mem['hF44D]=8'hF1; mem['hF44E]=8'h5E; mem['hF44F]=8'hD7;
    mem['hF450]=8'h50; mem['hF451]=8'hD7; mem['hF452]=8'h51; mem['hF453]=8'hD7;
    mem['hF454]=8'h52; mem['hF455]=8'hD7; mem['hF456]=8'h53; mem['hF457]=8'h39;
    mem['hF458]=8'h9E; mem['hF459]=8'h74; mem['hF45A]=8'h9F; mem['hF45B]=8'h54;
    mem['hF45C]=8'h9F; mem['hF45D]=8'h4F; mem['hF45E]=8'h9F; mem['hF45F]=8'h51;
    mem['hF460]=8'h9F; mem['hF461]=8'h52; mem['hF462]=8'h9F; mem['hF463]=8'h47;
    mem['hF464]=8'h9F; mem['hF465]=8'h45; mem['hF466]=8'h25; mem['hF467]=8'h64;
    mem['hF468]=8'hBD; mem['hF469]=8'hFB; mem['hF46A]=8'h95; mem['hF46B]=8'h81;
    mem['hF46C]=8'h2D; mem['hF46D]=8'h26; mem['hF46E]=8'h04; mem['hF46F]=8'h03;
    mem['hF470]=8'h55; mem['hF471]=8'h20; mem['hF472]=8'h04; mem['hF473]=8'h81;
    mem['hF474]=8'h2B; mem['hF475]=8'h26; mem['hF476]=8'h04; mem['hF477]=8'h9D;
    mem['hF478]=8'h7C; mem['hF479]=8'h25; mem['hF47A]=8'h51; mem['hF47B]=8'h81;
    mem['hF47C]=8'h2E; mem['hF47D]=8'h27; mem['hF47E]=8'h28; mem['hF47F]=8'h81;
    mem['hF480]=8'h45; mem['hF481]=8'h26; mem['hF482]=8'h28; mem['hF483]=8'h9D;
    mem['hF484]=8'h7C; mem['hF485]=8'h25; mem['hF486]=8'h64; mem['hF487]=8'h81;
    mem['hF488]=8'hA7; mem['hF489]=8'h27; mem['hF48A]=8'h0E; mem['hF48B]=8'h81;
    mem['hF48C]=8'h2D; mem['hF48D]=8'h27; mem['hF48E]=8'h0A; mem['hF48F]=8'h81;
    mem['hF490]=8'hA6; mem['hF491]=8'h27; mem['hF492]=8'h08; mem['hF493]=8'h81;
    mem['hF494]=8'h2B; mem['hF495]=8'h27; mem['hF496]=8'h04; mem['hF497]=8'h20;
    mem['hF498]=8'h06; mem['hF499]=8'h03; mem['hF49A]=8'h48; mem['hF49B]=8'h9D;
    mem['hF49C]=8'h7C; mem['hF49D]=8'h25; mem['hF49E]=8'h4C; mem['hF49F]=8'h0D;
    mem['hF4A0]=8'h48; mem['hF4A1]=8'h27; mem['hF4A2]=8'h08; mem['hF4A3]=8'h00;
    mem['hF4A4]=8'h47; mem['hF4A5]=8'h20; mem['hF4A6]=8'h04; mem['hF4A7]=8'h03;
    mem['hF4A8]=8'h46; mem['hF4A9]=8'h26; mem['hF4AA]=8'hCC; mem['hF4AB]=8'h96;
    mem['hF4AC]=8'h47; mem['hF4AD]=8'h90; mem['hF4AE]=8'h45; mem['hF4AF]=8'h97;
    mem['hF4B0]=8'h47; mem['hF4B1]=8'h27; mem['hF4B2]=8'h12; mem['hF4B3]=8'h2A;
    mem['hF4B4]=8'h09; mem['hF4B5]=8'hBD; mem['hF4B6]=8'hF2; mem['hF4B7]=8'hC8;
    mem['hF4B8]=8'h0C; mem['hF4B9]=8'h47; mem['hF4BA]=8'h26; mem['hF4BB]=8'hF9;
    mem['hF4BC]=8'h20; mem['hF4BD]=8'h07; mem['hF4BE]=8'hBD; mem['hF4BF]=8'hF2;
    mem['hF4C0]=8'hB0; mem['hF4C1]=8'h0A; mem['hF4C2]=8'h47; mem['hF4C3]=8'h26;
    mem['hF4C4]=8'hF9; mem['hF4C5]=8'h96; mem['hF4C6]=8'h55; mem['hF4C7]=8'h2A;
    mem['hF4C8]=8'h8E; mem['hF4C9]=8'h7E; mem['hF4CA]=8'hF6; mem['hF4CB]=8'h2F;
    mem['hF4CC]=8'hD6; mem['hF4CD]=8'h45; mem['hF4CE]=8'hD0; mem['hF4CF]=8'h46;
    mem['hF4D0]=8'hD7; mem['hF4D1]=8'h45; mem['hF4D2]=8'h34; mem['hF4D3]=8'h02;
    mem['hF4D4]=8'hBD; mem['hF4D5]=8'hF2; mem['hF4D6]=8'hB0; mem['hF4D7]=8'h35;
    mem['hF4D8]=8'h04; mem['hF4D9]=8'hC0; mem['hF4DA]=8'h30; mem['hF4DB]=8'h8D;
    mem['hF4DC]=8'h02; mem['hF4DD]=8'h20; mem['hF4DE]=8'h98; mem['hF4DF]=8'hBD;
    mem['hF4E0]=8'hF3; mem['hF4E1]=8'h75; mem['hF4E2]=8'hBD; mem['hF4E3]=8'hF3;
    mem['hF4E4]=8'hC2; mem['hF4E5]=8'h8E; mem['hF4E6]=8'h00; mem['hF4E7]=8'h40;
    mem['hF4E8]=8'h7E; mem['hF4E9]=8'hF1; mem['hF4EA]=8'h08; mem['hF4EB]=8'hD6;
    mem['hF4EC]=8'h47; mem['hF4ED]=8'h58; mem['hF4EE]=8'h58; mem['hF4EF]=8'hDB;
    mem['hF4F0]=8'h47; mem['hF4F1]=8'h58; mem['hF4F2]=8'h80; mem['hF4F3]=8'h30;
    mem['hF4F4]=8'h34; mem['hF4F5]=8'h04; mem['hF4F6]=8'hAB; mem['hF4F7]=8'hE0;
    mem['hF4F8]=8'h97; mem['hF4F9]=8'h47; mem['hF4FA]=8'h20; mem['hF4FB]=8'h9F;
    mem['hF4FC]=8'h9B; mem['hF4FD]=8'h3E; mem['hF4FE]=8'hBC; mem['hF4FF]=8'h1F;
    mem['hF500]=8'hFD; mem['hF501]=8'h9E; mem['hF502]=8'h6E; mem['hF503]=8'h6B;
    mem['hF504]=8'h27; mem['hF505]=8'hFD; mem['hF506]=8'h9E; mem['hF507]=8'h6E;
    mem['hF508]=8'h6B; mem['hF509]=8'h28; mem['hF50A]=8'h00; mem['hF50B]=8'h8E;
    mem['hF50C]=8'hE3; mem['hF50D]=8'hA4; mem['hF50E]=8'h8D; mem['hF50F]=8'h0C;
    mem['hF510]=8'hDC; mem['hF511]=8'h68; mem['hF512]=8'hDD; mem['hF513]=8'h50;
    mem['hF514]=8'hC6; mem['hF515]=8'h90; mem['hF516]=8'h43; mem['hF517]=8'hBD;
    mem['hF518]=8'hF3; mem['hF519]=8'hCC; mem['hF51A]=8'h8D; mem['hF51B]=8'h03;
    mem['hF51C]=8'h7E; mem['hF51D]=8'hF0; mem['hF51E]=8'hE2; mem['hF51F]=8'hCE;
    mem['hF520]=8'h01; mem['hF521]=8'hF1; mem['hF522]=8'h86; mem['hF523]=8'h20;
    mem['hF524]=8'hD6; mem['hF525]=8'h54; mem['hF526]=8'h2A; mem['hF527]=8'h02;
    mem['hF528]=8'h86; mem['hF529]=8'h2D; mem['hF52A]=8'hA7; mem['hF52B]=8'hC0;
    mem['hF52C]=8'hDF; mem['hF52D]=8'h64; mem['hF52E]=8'h97; mem['hF52F]=8'h54;
    mem['hF530]=8'h86; mem['hF531]=8'h30; mem['hF532]=8'hD6; mem['hF533]=8'h4F;
    mem['hF534]=8'h10; mem['hF535]=8'h27; mem['hF536]=8'h00; mem['hF537]=8'hC6;
    mem['hF538]=8'h4F; mem['hF539]=8'hC1; mem['hF53A]=8'h80; mem['hF53B]=8'h22;
    mem['hF53C]=8'h08; mem['hF53D]=8'h8E; mem['hF53E]=8'hF5; mem['hF53F]=8'h06;
    mem['hF540]=8'hBD; mem['hF541]=8'hF2; mem['hF542]=8'h10; mem['hF543]=8'h86;
    mem['hF544]=8'hF7; mem['hF545]=8'h97; mem['hF546]=8'h45; mem['hF547]=8'h8E;
    mem['hF548]=8'hF5; mem['hF549]=8'h01; mem['hF54A]=8'hBD; mem['hF54B]=8'hF3;
    mem['hF54C]=8'hE6; mem['hF54D]=8'h2E; mem['hF54E]=8'h0F; mem['hF54F]=8'h8E;
    mem['hF550]=8'hF4; mem['hF551]=8'hFC; mem['hF552]=8'hBD; mem['hF553]=8'hF3;
    mem['hF554]=8'hE6; mem['hF555]=8'h2E; mem['hF556]=8'h0E; mem['hF557]=8'hBD;
    mem['hF558]=8'hF2; mem['hF559]=8'hB0; mem['hF55A]=8'h0A; mem['hF55B]=8'h45;
    mem['hF55C]=8'h20; mem['hF55D]=8'hF1; mem['hF55E]=8'hBD; mem['hF55F]=8'hF2;
    mem['hF560]=8'hC8; mem['hF561]=8'h0C; mem['hF562]=8'h45; mem['hF563]=8'h20;
    mem['hF564]=8'hE2; mem['hF565]=8'hBD; mem['hF566]=8'hF0; mem['hF567]=8'hFA;
    mem['hF568]=8'hBD; mem['hF569]=8'hF4; mem['hF56A]=8'h0E; mem['hF56B]=8'hC6;
    mem['hF56C]=8'h01; mem['hF56D]=8'h96; mem['hF56E]=8'h45; mem['hF56F]=8'h8B;
    mem['hF570]=8'h0A; mem['hF571]=8'h2B; mem['hF572]=8'h09; mem['hF573]=8'h81;
    mem['hF574]=8'h0B; mem['hF575]=8'h24; mem['hF576]=8'h05; mem['hF577]=8'h4A;
    mem['hF578]=8'h1F; mem['hF579]=8'h89; mem['hF57A]=8'h86; mem['hF57B]=8'h02;
    mem['hF57C]=8'h4A; mem['hF57D]=8'h4A; mem['hF57E]=8'h97; mem['hF57F]=8'h47;
    mem['hF580]=8'hD7; mem['hF581]=8'h45; mem['hF582]=8'h2E; mem['hF583]=8'h0D;
    mem['hF584]=8'hDE; mem['hF585]=8'h64; mem['hF586]=8'h86; mem['hF587]=8'h2E;
    mem['hF588]=8'hA7; mem['hF589]=8'hC0; mem['hF58A]=8'h5D; mem['hF58B]=8'h27;
    mem['hF58C]=8'h04; mem['hF58D]=8'h86; mem['hF58E]=8'h30; mem['hF58F]=8'hA7;
    mem['hF590]=8'hC0; mem['hF591]=8'h8E; mem['hF592]=8'hF6; mem['hF593]=8'h0B;
    mem['hF594]=8'hC6; mem['hF595]=8'h80; mem['hF596]=8'h96; mem['hF597]=8'h53;
    mem['hF598]=8'hAB; mem['hF599]=8'h03; mem['hF59A]=8'h97; mem['hF59B]=8'h53;
    mem['hF59C]=8'h96; mem['hF59D]=8'h52; mem['hF59E]=8'hA9; mem['hF59F]=8'h02;
    mem['hF5A0]=8'h97; mem['hF5A1]=8'h52; mem['hF5A2]=8'h96; mem['hF5A3]=8'h51;
    mem['hF5A4]=8'hA9; mem['hF5A5]=8'h01; mem['hF5A6]=8'h97; mem['hF5A7]=8'h51;
    mem['hF5A8]=8'h96; mem['hF5A9]=8'h50; mem['hF5AA]=8'hA9; mem['hF5AB]=8'h84;
    mem['hF5AC]=8'h97; mem['hF5AD]=8'h50; mem['hF5AE]=8'h5C; mem['hF5AF]=8'h56;
    mem['hF5B0]=8'h59; mem['hF5B1]=8'h28; mem['hF5B2]=8'hE3; mem['hF5B3]=8'h24;
    mem['hF5B4]=8'h03; mem['hF5B5]=8'hC0; mem['hF5B6]=8'h0B; mem['hF5B7]=8'h50;
    mem['hF5B8]=8'hCB; mem['hF5B9]=8'h2F; mem['hF5BA]=8'h30; mem['hF5BB]=8'h04;
    mem['hF5BC]=8'h1F; mem['hF5BD]=8'h98; mem['hF5BE]=8'h84; mem['hF5BF]=8'h7F;
    mem['hF5C0]=8'hA7; mem['hF5C1]=8'hC0; mem['hF5C2]=8'h0A; mem['hF5C3]=8'h45;
    mem['hF5C4]=8'h26; mem['hF5C5]=8'h04; mem['hF5C6]=8'h86; mem['hF5C7]=8'h2E;
    mem['hF5C8]=8'hA7; mem['hF5C9]=8'hC0; mem['hF5CA]=8'h53; mem['hF5CB]=8'hC4;
    mem['hF5CC]=8'h80; mem['hF5CD]=8'h8C; mem['hF5CE]=8'hF6; mem['hF5CF]=8'h2F;
    mem['hF5D0]=8'h26; mem['hF5D1]=8'hC4; mem['hF5D2]=8'hA6; mem['hF5D3]=8'hC2;
    mem['hF5D4]=8'h81; mem['hF5D5]=8'h30; mem['hF5D6]=8'h27; mem['hF5D7]=8'hFA;
    mem['hF5D8]=8'h81; mem['hF5D9]=8'h2E; mem['hF5DA]=8'h26; mem['hF5DB]=8'h02;
    mem['hF5DC]=8'h33; mem['hF5DD]=8'h5F; mem['hF5DE]=8'h86; mem['hF5DF]=8'h2B;
    mem['hF5E0]=8'hD6; mem['hF5E1]=8'h47; mem['hF5E2]=8'h27; mem['hF5E3]=8'h1C;
    mem['hF5E4]=8'h2A; mem['hF5E5]=8'h03; mem['hF5E6]=8'h86; mem['hF5E7]=8'h2D;
    mem['hF5E8]=8'h50; mem['hF5E9]=8'hA7; mem['hF5EA]=8'h42; mem['hF5EB]=8'h86;
    mem['hF5EC]=8'h45; mem['hF5ED]=8'hA7; mem['hF5EE]=8'h41; mem['hF5EF]=8'h86;
    mem['hF5F0]=8'h2F; mem['hF5F1]=8'h4C; mem['hF5F2]=8'hC0; mem['hF5F3]=8'h0A;
    mem['hF5F4]=8'h24; mem['hF5F5]=8'hFB; mem['hF5F6]=8'hCB; mem['hF5F7]=8'h3A;
    mem['hF5F8]=8'hED; mem['hF5F9]=8'h43; mem['hF5FA]=8'h6F; mem['hF5FB]=8'h45;
    mem['hF5FC]=8'h20; mem['hF5FD]=8'h04; mem['hF5FE]=8'hA7; mem['hF5FF]=8'hC4;
    mem['hF600]=8'h6F; mem['hF601]=8'h41; mem['hF602]=8'h8E; mem['hF603]=8'h01;
    mem['hF604]=8'hF1; mem['hF605]=8'h39; mem['hF606]=8'h80; mem['hF607]=8'h00;
    mem['hF608]=8'h00; mem['hF609]=8'h00; mem['hF60A]=8'h00; mem['hF60B]=8'hFA;
    mem['hF60C]=8'h0A; mem['hF60D]=8'h1F; mem['hF60E]=8'h00; mem['hF60F]=8'h00;
    mem['hF610]=8'h98; mem['hF611]=8'h96; mem['hF612]=8'h80; mem['hF613]=8'hFF;
    mem['hF614]=8'hF0; mem['hF615]=8'hBD; mem['hF616]=8'hC0; mem['hF617]=8'h00;
    mem['hF618]=8'h01; mem['hF619]=8'h86; mem['hF61A]=8'hA0; mem['hF61B]=8'hFF;
    mem['hF61C]=8'hFF; mem['hF61D]=8'hD8; mem['hF61E]=8'hF0; mem['hF61F]=8'h00;
    mem['hF620]=8'h00; mem['hF621]=8'h03; mem['hF622]=8'hE8; mem['hF623]=8'hFF;
    mem['hF624]=8'hFF; mem['hF625]=8'hFF; mem['hF626]=8'h9C; mem['hF627]=8'h00;
    mem['hF628]=8'h00; mem['hF629]=8'h00; mem['hF62A]=8'h0A; mem['hF62B]=8'hFF;
    mem['hF62C]=8'hFF; mem['hF62D]=8'hFF; mem['hF62E]=8'hFF; mem['hF62F]=8'h96;
    mem['hF630]=8'h4F; mem['hF631]=8'h27; mem['hF632]=8'h02; mem['hF633]=8'h03;
    mem['hF634]=8'h54; mem['hF635]=8'h39; mem['hF636]=8'h9F; mem['hF637]=8'h64;
    mem['hF638]=8'hBD; mem['hF639]=8'hF3; mem['hF63A]=8'h75; mem['hF63B]=8'h8D;
    mem['hF63C]=8'h05; mem['hF63D]=8'h8D; mem['hF63E]=8'h08; mem['hF63F]=8'h8E;
    mem['hF640]=8'h00; mem['hF641]=8'h40; mem['hF642]=8'h7E; mem['hF643]=8'hF2;
    mem['hF644]=8'h10; mem['hF645]=8'h9F; mem['hF646]=8'h64; mem['hF647]=8'hBD;
    mem['hF648]=8'hF3; mem['hF649]=8'h70; mem['hF64A]=8'h9E; mem['hF64B]=8'h64;
    mem['hF64C]=8'hE6; mem['hF64D]=8'h80; mem['hF64E]=8'hD7; mem['hF64F]=8'h55;
    mem['hF650]=8'h9F; mem['hF651]=8'h64; mem['hF652]=8'h8D; mem['hF653]=8'hEE;
    mem['hF654]=8'h9E; mem['hF655]=8'h64; mem['hF656]=8'h30; mem['hF657]=8'h05;
    mem['hF658]=8'h9F; mem['hF659]=8'h64; mem['hF65A]=8'hBD; mem['hF65B]=8'hF1;
    mem['hF65C]=8'h08; mem['hF65D]=8'h8E; mem['hF65E]=8'h00; mem['hF65F]=8'h45;
    mem['hF660]=8'h0A; mem['hF661]=8'h55; mem['hF662]=8'h26; mem['hF663]=8'hEE;
    mem['hF664]=8'h39; mem['hF665]=8'hBD; mem['hF666]=8'hF3; mem['hF667]=8'hB3;
    mem['hF668]=8'h2B; mem['hF669]=8'h1F; mem['hF66A]=8'h27; mem['hF66B]=8'h15;
    mem['hF66C]=8'h8D; mem['hF66D]=8'h10; mem['hF66E]=8'hBD; mem['hF66F]=8'hF3;
    mem['hF670]=8'h75; mem['hF671]=8'h8D; mem['hF672]=8'h0E; mem['hF673]=8'h8E;
    mem['hF674]=8'h00; mem['hF675]=8'h40; mem['hF676]=8'h8D; mem['hF677]=8'hCA;
    mem['hF678]=8'h8E; mem['hF679]=8'hF2; mem['hF67A]=8'h0B; mem['hF67B]=8'hBD;
    mem['hF67C]=8'hF1; mem['hF67D]=8'h08; mem['hF67E]=8'h7E; mem['hF67F]=8'hF4;
    mem['hF680]=8'h34; mem['hF681]=8'h9E; mem['hF682]=8'hB1; mem['hF683]=8'h9F;
    mem['hF684]=8'h50; mem['hF685]=8'h9E; mem['hF686]=8'hB3; mem['hF687]=8'h9F;
    mem['hF688]=8'h52; mem['hF689]=8'hBE; mem['hF68A]=8'hF6; mem['hF68B]=8'hB6;
    mem['hF68C]=8'h9F; mem['hF68D]=8'h5D; mem['hF68E]=8'hBE; mem['hF68F]=8'hF6;
    mem['hF690]=8'hB8; mem['hF691]=8'h9F; mem['hF692]=8'h5F; mem['hF693]=8'hBD;
    mem['hF694]=8'hF2; mem['hF695]=8'h16; mem['hF696]=8'hDC; mem['hF697]=8'h8A;
    mem['hF698]=8'hC3; mem['hF699]=8'h65; mem['hF69A]=8'h8B; mem['hF69B]=8'hDD;
    mem['hF69C]=8'hB3; mem['hF69D]=8'hDD; mem['hF69E]=8'h52; mem['hF69F]=8'hDC;
    mem['hF6A0]=8'h88; mem['hF6A1]=8'hC9; mem['hF6A2]=8'hB0; mem['hF6A3]=8'h89;
    mem['hF6A4]=8'h05; mem['hF6A5]=8'hDD; mem['hF6A6]=8'hB1; mem['hF6A7]=8'hDD;
    mem['hF6A8]=8'h50; mem['hF6A9]=8'h0F; mem['hF6AA]=8'h54; mem['hF6AB]=8'h86;
    mem['hF6AC]=8'h80; mem['hF6AD]=8'h97; mem['hF6AE]=8'h4F; mem['hF6AF]=8'h96;
    mem['hF6B0]=8'h15; mem['hF6B1]=8'h97; mem['hF6B2]=8'h63; mem['hF6B3]=8'h7E;
    mem['hF6B4]=8'hF1; mem['hF6B5]=8'h62; mem['hF6B6]=8'h40; mem['hF6B7]=8'hE6;
    mem['hF6B8]=8'h4D; mem['hF6B9]=8'hAB; mem['hF6BA]=8'hBD; mem['hF6BB]=8'hF3;
    mem['hF6BC]=8'hA5; mem['hF6BD]=8'h8E; mem['hF6BE]=8'hF6; mem['hF6BF]=8'hFF;
    mem['hF6C0]=8'hD6; mem['hF6C1]=8'h61; mem['hF6C2]=8'hBD; mem['hF6C3]=8'hF2;
    mem['hF6C4]=8'hCF; mem['hF6C5]=8'hBD; mem['hF6C6]=8'hF3; mem['hF6C7]=8'hA5;
    mem['hF6C8]=8'h8D; mem['hF6C9]=8'hB4; mem['hF6CA]=8'h0F; mem['hF6CB]=8'h62;
    mem['hF6CC]=8'h96; mem['hF6CD]=8'h5C; mem['hF6CE]=8'hD6; mem['hF6CF]=8'h4F;
    mem['hF6D0]=8'hBD; mem['hF6D1]=8'hF1; mem['hF6D2]=8'h02; mem['hF6D3]=8'h8E;
    mem['hF6D4]=8'hF7; mem['hF6D5]=8'h04; mem['hF6D6]=8'hBD; mem['hF6D7]=8'hF0;
    mem['hF6D8]=8'hFF; mem['hF6D9]=8'h96; mem['hF6DA]=8'h54; mem['hF6DB]=8'h34;
    mem['hF6DC]=8'h02; mem['hF6DD]=8'h2A; mem['hF6DE]=8'h09; mem['hF6DF]=8'hBD;
    mem['hF6E0]=8'hF0; mem['hF6E1]=8'hFA; mem['hF6E2]=8'h96; mem['hF6E3]=8'h54;
    mem['hF6E4]=8'h2B; mem['hF6E5]=8'h05; mem['hF6E6]=8'h03; mem['hF6E7]=8'h0A;
    mem['hF6E8]=8'hBD; mem['hF6E9]=8'hF6; mem['hF6EA]=8'h2F; mem['hF6EB]=8'h8E;
    mem['hF6EC]=8'hF7; mem['hF6ED]=8'h04; mem['hF6EE]=8'hBD; mem['hF6EF]=8'hF1;
    mem['hF6F0]=8'h08; mem['hF6F1]=8'h35; mem['hF6F2]=8'h02; mem['hF6F3]=8'h4D;
    mem['hF6F4]=8'h2A; mem['hF6F5]=8'h03; mem['hF6F6]=8'hBD; mem['hF6F7]=8'hF6;
    mem['hF6F8]=8'h2F; mem['hF6F9]=8'h8E; mem['hF6FA]=8'hF7; mem['hF6FB]=8'h09;
    mem['hF6FC]=8'h7E; mem['hF6FD]=8'hF6; mem['hF6FE]=8'h36; mem['hF6FF]=8'h83;
    mem['hF700]=8'h49; mem['hF701]=8'h0F; mem['hF702]=8'hDA; mem['hF703]=8'hA2;
    mem['hF704]=8'h7F; mem['hF705]=8'h00; mem['hF706]=8'h00; mem['hF707]=8'h00;
    mem['hF708]=8'h00; mem['hF709]=8'h05; mem['hF70A]=8'h84; mem['hF70B]=8'hE6;
    mem['hF70C]=8'h1A; mem['hF70D]=8'h2D; mem['hF70E]=8'h1B; mem['hF70F]=8'h86;
    mem['hF710]=8'h28; mem['hF711]=8'h07; mem['hF712]=8'hFB; mem['hF713]=8'hF8;
    mem['hF714]=8'h87; mem['hF715]=8'h99; mem['hF716]=8'h68; mem['hF717]=8'h89;
    mem['hF718]=8'h01; mem['hF719]=8'h87; mem['hF71A]=8'h23; mem['hF71B]=8'h35;
    mem['hF71C]=8'hDF; mem['hF71D]=8'hE1; mem['hF71E]=8'h86; mem['hF71F]=8'hA5;
    mem['hF720]=8'h5D; mem['hF721]=8'hE7; mem['hF722]=8'h28; mem['hF723]=8'h83;
    mem['hF724]=8'h49; mem['hF725]=8'h0F; mem['hF726]=8'hDA; mem['hF727]=8'hA2;
    mem['hF728]=8'hA1; mem['hF729]=8'h54; mem['hF72A]=8'h46; mem['hF72B]=8'h8F;
    mem['hF72C]=8'h13; mem['hF72D]=8'h8F; mem['hF72E]=8'h52; mem['hF72F]=8'h43;
    mem['hF730]=8'h89; mem['hF731]=8'hCD; mem['hF732]=8'h8E; mem['hF733]=8'hF7;
    mem['hF734]=8'h65; mem['hF735]=8'hBD; mem['hF736]=8'hF1; mem['hF737]=8'h08;
    mem['hF738]=8'h7E; mem['hF739]=8'hF6; mem['hF73A]=8'hBA; mem['hF73B]=8'hBD;
    mem['hF73C]=8'hF3; mem['hF73D]=8'h75; mem['hF73E]=8'h0F; mem['hF73F]=8'h0A;
    mem['hF740]=8'h8D; mem['hF741]=8'hF6; mem['hF742]=8'h8E; mem['hF743]=8'h00;
    mem['hF744]=8'h4A; mem['hF745]=8'hBD; mem['hF746]=8'hF3; mem['hF747]=8'h7B;
    mem['hF748]=8'h8E; mem['hF749]=8'h00; mem['hF74A]=8'h40; mem['hF74B]=8'hBD;
    mem['hF74C]=8'hF3; mem['hF74D]=8'h5A; mem['hF74E]=8'h0F; mem['hF74F]=8'h54;
    mem['hF750]=8'h96; mem['hF751]=8'h0A; mem['hF752]=8'h8D; mem['hF753]=8'h0C;
    mem['hF754]=8'h0D; mem['hF755]=8'h4F; mem['hF756]=8'h10; mem['hF757]=8'h27;
    mem['hF758]=8'hFA; mem['hF759]=8'h7E; mem['hF75A]=8'h8E; mem['hF75B]=8'h00;
    mem['hF75C]=8'h4A; mem['hF75D]=8'h7E; mem['hF75E]=8'hF2; mem['hF75F]=8'hD5;
    mem['hF760]=8'h34; mem['hF761]=8'h02; mem['hF762]=8'h7E; mem['hF763]=8'hF6;
    mem['hF764]=8'hE8; mem['hF765]=8'h81; mem['hF766]=8'h49; mem['hF767]=8'h0F;
    mem['hF768]=8'hDA; mem['hF769]=8'hA2; mem['hF76A]=8'h96; mem['hF76B]=8'h54;
    mem['hF76C]=8'h34; mem['hF76D]=8'h02; mem['hF76E]=8'h2A; mem['hF76F]=8'h02;
    mem['hF770]=8'h8D; mem['hF771]=8'h24; mem['hF772]=8'h96; mem['hF773]=8'h4F;
    mem['hF774]=8'h34; mem['hF775]=8'h02; mem['hF776]=8'h81; mem['hF777]=8'h81;
    mem['hF778]=8'h25; mem['hF779]=8'h05; mem['hF77A]=8'h8E; mem['hF77B]=8'hF2;
    mem['hF77C]=8'h0B; mem['hF77D]=8'h8D; mem['hF77E]=8'hDE; mem['hF77F]=8'h8E;
    mem['hF780]=8'hF7; mem['hF781]=8'h9A; mem['hF782]=8'hBD; mem['hF783]=8'hF6;
    mem['hF784]=8'h36; mem['hF785]=8'h35; mem['hF786]=8'h02; mem['hF787]=8'h81;
    mem['hF788]=8'h81; mem['hF789]=8'h25; mem['hF78A]=8'h06; mem['hF78B]=8'h8E;
    mem['hF78C]=8'hF7; mem['hF78D]=8'h65; mem['hF78E]=8'hBD; mem['hF78F]=8'hF0;
    mem['hF790]=8'hFF; mem['hF791]=8'h35; mem['hF792]=8'h02; mem['hF793]=8'h4D;
    mem['hF794]=8'h2A; mem['hF795]=8'h03; mem['hF796]=8'h7E; mem['hF797]=8'hF6;
    mem['hF798]=8'h2F; mem['hF799]=8'h39; mem['hF79A]=8'h0B; mem['hF79B]=8'h76;
    mem['hF79C]=8'hB3; mem['hF79D]=8'h83; mem['hF79E]=8'hBD; mem['hF79F]=8'hD3;
    mem['hF7A0]=8'h79; mem['hF7A1]=8'h1E; mem['hF7A2]=8'hF4; mem['hF7A3]=8'hA6;
    mem['hF7A4]=8'hF5; mem['hF7A5]=8'h7B; mem['hF7A6]=8'h83; mem['hF7A7]=8'hFC;
    mem['hF7A8]=8'hB0; mem['hF7A9]=8'h10; mem['hF7AA]=8'h7C; mem['hF7AB]=8'h0C;
    mem['hF7AC]=8'h1F; mem['hF7AD]=8'h67; mem['hF7AE]=8'hCA; mem['hF7AF]=8'h7C;
    mem['hF7B0]=8'hDE; mem['hF7B1]=8'h53; mem['hF7B2]=8'hCB; mem['hF7B3]=8'hC1;
    mem['hF7B4]=8'h7D; mem['hF7B5]=8'h14; mem['hF7B6]=8'h64; mem['hF7B7]=8'h70;
    mem['hF7B8]=8'h4C; mem['hF7B9]=8'h7D; mem['hF7BA]=8'hB7; mem['hF7BB]=8'hEA;
    mem['hF7BC]=8'h51; mem['hF7BD]=8'h7A; mem['hF7BE]=8'h7D; mem['hF7BF]=8'h63;
    mem['hF7C0]=8'h30; mem['hF7C1]=8'h88; mem['hF7C2]=8'h7E; mem['hF7C3]=8'h7E;
    mem['hF7C4]=8'h92; mem['hF7C5]=8'h44; mem['hF7C6]=8'h99; mem['hF7C7]=8'h3A;
    mem['hF7C8]=8'h7E; mem['hF7C9]=8'h4C; mem['hF7CA]=8'hCC; mem['hF7CB]=8'h91;
    mem['hF7CC]=8'hC7; mem['hF7CD]=8'h7F; mem['hF7CE]=8'hAA; mem['hF7CF]=8'hAA;
    mem['hF7D0]=8'hAA; mem['hF7D1]=8'h13; mem['hF7D2]=8'h81; mem['hF7D3]=8'h00;
    mem['hF7D4]=8'h00; mem['hF7D5]=8'h00; mem['hF7D6]=8'h00; mem['hF7D7]=8'h03;
    mem['hF7D8]=8'h7F; mem['hF7D9]=8'h5E; mem['hF7DA]=8'h56; mem['hF7DB]=8'hCB;
    mem['hF7DC]=8'h79; mem['hF7DD]=8'h80; mem['hF7DE]=8'h13; mem['hF7DF]=8'h9B;
    mem['hF7E0]=8'h0B; mem['hF7E1]=8'h64; mem['hF7E2]=8'h80; mem['hF7E3]=8'h76;
    mem['hF7E4]=8'h38; mem['hF7E5]=8'h93; mem['hF7E6]=8'h16; mem['hF7E7]=8'h82;
    mem['hF7E8]=8'h38; mem['hF7E9]=8'hAA; mem['hF7EA]=8'h3B; mem['hF7EB]=8'h20;
    mem['hF7EC]=8'h80; mem['hF7ED]=8'h35; mem['hF7EE]=8'h04; mem['hF7EF]=8'hF3;
    mem['hF7F0]=8'h34; mem['hF7F1]=8'h81; mem['hF7F2]=8'h35; mem['hF7F3]=8'h04;
    mem['hF7F4]=8'hF3; mem['hF7F5]=8'h34; mem['hF7F6]=8'h80; mem['hF7F7]=8'h80;
    mem['hF7F8]=8'h00; mem['hF7F9]=8'h00; mem['hF7FA]=8'h00; mem['hF7FB]=8'h80;
    mem['hF7FC]=8'h31; mem['hF7FD]=8'h72; mem['hF7FE]=8'h17; mem['hF7FF]=8'hF8;
    mem['hF800]=8'hBD; mem['hF801]=8'hF3; mem['hF802]=8'hB3; mem['hF803]=8'h10;
    mem['hF804]=8'h2F; mem['hF805]=8'hF3; mem['hF806]=8'hC7; mem['hF807]=8'h8E;
    mem['hF808]=8'hF7; mem['hF809]=8'hEC; mem['hF80A]=8'h96; mem['hF80B]=8'h4F;
    mem['hF80C]=8'h80; mem['hF80D]=8'h80; mem['hF80E]=8'h34; mem['hF80F]=8'h02;
    mem['hF810]=8'h86; mem['hF811]=8'h80; mem['hF812]=8'h97; mem['hF813]=8'h4F;
    mem['hF814]=8'hBD; mem['hF815]=8'hF1; mem['hF816]=8'h08; mem['hF817]=8'h8E;
    mem['hF818]=8'hF7; mem['hF819]=8'hF1; mem['hF81A]=8'hBD; mem['hF81B]=8'hF2;
    mem['hF81C]=8'hD5; mem['hF81D]=8'h8E; mem['hF81E]=8'hF2; mem['hF81F]=8'h0B;
    mem['hF820]=8'hBD; mem['hF821]=8'hF0; mem['hF822]=8'hFF; mem['hF823]=8'h8E;
    mem['hF824]=8'hF7; mem['hF825]=8'hD7; mem['hF826]=8'hBD; mem['hF827]=8'hF6;
    mem['hF828]=8'h36; mem['hF829]=8'h8E; mem['hF82A]=8'hF7; mem['hF82B]=8'hF6;
    mem['hF82C]=8'hBD; mem['hF82D]=8'hF1; mem['hF82E]=8'h08; mem['hF82F]=8'h35;
    mem['hF830]=8'h04; mem['hF831]=8'hBD; mem['hF832]=8'hF4; mem['hF833]=8'hDF;
    mem['hF834]=8'h8E; mem['hF835]=8'hF7; mem['hF836]=8'hFB; mem['hF837]=8'h7E;
    mem['hF838]=8'hF2; mem['hF839]=8'h10; mem['hF83A]=8'hBD; mem['hF83B]=8'hF3;
    mem['hF83C]=8'hA5; mem['hF83D]=8'h8E; mem['hF83E]=8'hF6; mem['hF83F]=8'h06;
    mem['hF840]=8'hBD; mem['hF841]=8'hF3; mem['hF842]=8'h5A; mem['hF843]=8'h27;
    mem['hF844]=8'h67; mem['hF845]=8'h4D; mem['hF846]=8'h26; mem['hF847]=8'h03;
    mem['hF848]=8'h7E; mem['hF849]=8'hF1; mem['hF84A]=8'h80; mem['hF84B]=8'h8E;
    mem['hF84C]=8'h00; mem['hF84D]=8'h4A; mem['hF84E]=8'hBD; mem['hF84F]=8'hF3;
    mem['hF850]=8'h7B; mem['hF851]=8'h5F; mem['hF852]=8'h96; mem['hF853]=8'h61;
    mem['hF854]=8'h2A; mem['hF855]=8'h10; mem['hF856]=8'hBD; mem['hF857]=8'hF4;
    mem['hF858]=8'h34; mem['hF859]=8'h8E; mem['hF85A]=8'h00; mem['hF85B]=8'h4A;
    mem['hF85C]=8'h96; mem['hF85D]=8'h61; mem['hF85E]=8'hBD; mem['hF85F]=8'hF3;
    mem['hF860]=8'hE6; mem['hF861]=8'h26; mem['hF862]=8'h03; mem['hF863]=8'h43;
    mem['hF864]=8'hD6; mem['hF865]=8'h01; mem['hF866]=8'hBD; mem['hF867]=8'hF3;
    mem['hF868]=8'h92; mem['hF869]=8'h34; mem['hF86A]=8'h04; mem['hF86B]=8'hBD;
    mem['hF86C]=8'hF8; mem['hF86D]=8'h00; mem['hF86E]=8'h8E; mem['hF86F]=8'h00;
    mem['hF870]=8'h4A; mem['hF871]=8'hBD; mem['hF872]=8'hF2; mem['hF873]=8'h10;
    mem['hF874]=8'h8D; mem['hF875]=8'h36; mem['hF876]=8'h35; mem['hF877]=8'h02;
    mem['hF878]=8'h46; mem['hF879]=8'h10; mem['hF87A]=8'h25; mem['hF87B]=8'hFD;
    mem['hF87C]=8'hB2; mem['hF87D]=8'h39; mem['hF87E]=8'h81; mem['hF87F]=8'h38;
    mem['hF880]=8'hAA; mem['hF881]=8'h3B; mem['hF882]=8'h29; mem['hF883]=8'h07;
    mem['hF884]=8'h71; mem['hF885]=8'h34; mem['hF886]=8'h58; mem['hF887]=8'h3E;
    mem['hF888]=8'h56; mem['hF889]=8'h74; mem['hF88A]=8'h16; mem['hF88B]=8'h7E;
    mem['hF88C]=8'hB3; mem['hF88D]=8'h1B; mem['hF88E]=8'h77; mem['hF88F]=8'h2F;
    mem['hF890]=8'hEE; mem['hF891]=8'hE3; mem['hF892]=8'h85; mem['hF893]=8'h7A;
    mem['hF894]=8'h1D; mem['hF895]=8'h84; mem['hF896]=8'h1C; mem['hF897]=8'h2A;
    mem['hF898]=8'h7C; mem['hF899]=8'h63; mem['hF89A]=8'h59; mem['hF89B]=8'h58;
    mem['hF89C]=8'h0A; mem['hF89D]=8'h7E; mem['hF89E]=8'h75; mem['hF89F]=8'hFD;
    mem['hF8A0]=8'hE7; mem['hF8A1]=8'hC6; mem['hF8A2]=8'h80; mem['hF8A3]=8'h31;
    mem['hF8A4]=8'h72; mem['hF8A5]=8'h18; mem['hF8A6]=8'h10; mem['hF8A7]=8'h81;
    mem['hF8A8]=8'h00; mem['hF8A9]=8'h00; mem['hF8AA]=8'h00; mem['hF8AB]=8'h00;
    mem['hF8AC]=8'h8E; mem['hF8AD]=8'hF8; mem['hF8AE]=8'h7E; mem['hF8AF]=8'hBD;
    mem['hF8B0]=8'hF2; mem['hF8B1]=8'h10; mem['hF8B2]=8'hBD; mem['hF8B3]=8'hF3;
    mem['hF8B4]=8'h75; mem['hF8B5]=8'h96; mem['hF8B6]=8'h4F; mem['hF8B7]=8'h81;
    mem['hF8B8]=8'h88; mem['hF8B9]=8'h25; mem['hF8BA]=8'h03; mem['hF8BB]=8'h7E;
    mem['hF8BC]=8'hF2; mem['hF8BD]=8'hA2; mem['hF8BE]=8'hBD; mem['hF8BF]=8'hF4;
    mem['hF8C0]=8'h34; mem['hF8C1]=8'h96; mem['hF8C2]=8'h01; mem['hF8C3]=8'h8B;
    mem['hF8C4]=8'h81; mem['hF8C5]=8'h27; mem['hF8C6]=8'hF4; mem['hF8C7]=8'h4A;
    mem['hF8C8]=8'h34; mem['hF8C9]=8'h02; mem['hF8CA]=8'h8E; mem['hF8CB]=8'h00;
    mem['hF8CC]=8'h40; mem['hF8CD]=8'hBD; mem['hF8CE]=8'hF0; mem['hF8CF]=8'hFF;
    mem['hF8D0]=8'h8E; mem['hF8D1]=8'hF8; mem['hF8D2]=8'h83; mem['hF8D3]=8'hBD;
    mem['hF8D4]=8'hF6; mem['hF8D5]=8'h45; mem['hF8D6]=8'h0F; mem['hF8D7]=8'h62;
    mem['hF8D8]=8'h35; mem['hF8D9]=8'h02; mem['hF8DA]=8'hBD; mem['hF8DB]=8'hF2;
    mem['hF8DC]=8'h8E; mem['hF8DD]=8'h39; mem['hF8DE]=8'hBD; mem['hF8DF]=8'hF3;
    mem['hF8E0]=8'hB3; mem['hF8E1]=8'h2B; mem['hF8E2]=8'h03; mem['hF8E3]=8'h7E;
    mem['hF8E4]=8'hF4; mem['hF8E5]=8'h34; mem['hF8E6]=8'h03; mem['hF8E7]=8'h54;
    mem['hF8E8]=8'h8D; mem['hF8E9]=8'hF9; mem['hF8EA]=8'h7E; mem['hF8EB]=8'hF6;
    mem['hF8EC]=8'h2F; mem['hF8ED]=8'hBD; mem['hF8EE]=8'hFD; mem['hF8EF]=8'h1B;
    mem['hF8F0]=8'h32; mem['hF8F1]=8'h62; mem['hF8F2]=8'h86; mem['hF8F3]=8'h01;
    mem['hF8F4]=8'h97; mem['hF8F5]=8'h98; mem['hF8F6]=8'hBD; mem['hF8F7]=8'hE4;
    mem['hF8F8]=8'hA2; mem['hF8F9]=8'h10; mem['hF8FA]=8'h25; mem['hF8FB]=8'hED;
    mem['hF8FC]=8'h82; mem['hF8FD]=8'hBD; mem['hF8FE]=8'hEF; mem['hF8FF]=8'h3B;
    mem['hF900]=8'h1F; mem['hF901]=8'h20; mem['hF902]=8'h83; mem['hF903]=8'h00;
    mem['hF904]=8'hF5; mem['hF905]=8'hD7; mem['hF906]=8'h97; mem['hF907]=8'hDC;
    mem['hF908]=8'h2B; mem['hF909]=8'hBD; mem['hF90A]=8'hF5; mem['hF90B]=8'h12;
    mem['hF90C]=8'hBD; mem['hF90D]=8'hF0; mem['hF90E]=8'hF2; mem['hF90F]=8'h8E;
    mem['hF910]=8'h00; mem['hF911]=8'hF4; mem['hF912]=8'hD6; mem['hF913]=8'h98;
    mem['hF914]=8'h26; mem['hF915]=8'h25; mem['hF916]=8'h5F; mem['hF917]=8'hBD;
    mem['hF918]=8'hFA; mem['hF919]=8'h41; mem['hF91A]=8'hBD; mem['hF91B]=8'hFF;
    mem['hF91C]=8'h73; mem['hF91D]=8'h25; mem['hF91E]=8'h0B; mem['hF91F]=8'h80;
    mem['hF920]=8'h30; mem['hF921]=8'h34; mem['hF922]=8'h02; mem['hF923]=8'h86;
    mem['hF924]=8'h0A; mem['hF925]=8'h3D; mem['hF926]=8'hEB; mem['hF927]=8'hE0;
    mem['hF928]=8'h20; mem['hF929]=8'hED; mem['hF92A]=8'hC0; mem['hF92B]=8'h01;
    mem['hF92C]=8'hC9; mem['hF92D]=8'h01; mem['hF92E]=8'h81; mem['hF92F]=8'h41;
    mem['hF930]=8'h26; mem['hF931]=8'h05; mem['hF932]=8'hBD; mem['hF933]=8'hF0;
    mem['hF934]=8'hA2; mem['hF935]=8'h20; mem['hF936]=8'hBB; mem['hF937]=8'h81;
    mem['hF938]=8'h4C; mem['hF939]=8'h26; mem['hF93A]=8'h0B; mem['hF93B]=8'h8D;
    mem['hF93C]=8'h31; mem['hF93D]=8'h0F; mem['hF93E]=8'h98; mem['hF93F]=8'hBD;
    mem['hF940]=8'hF0; mem['hF941]=8'hA2; mem['hF942]=8'h20; mem['hF943]=8'hC3;
    mem['hF944]=8'h32; mem['hF945]=8'h62; mem['hF946]=8'h81; mem['hF947]=8'h0D;
    mem['hF948]=8'h26; mem['hF949]=8'h0D; mem['hF94A]=8'h8D; mem['hF94B]=8'h22;
    mem['hF94C]=8'hBD; mem['hF94D]=8'hF0; mem['hF94E]=8'hA2; mem['hF94F]=8'h8E;
    mem['hF950]=8'h00; mem['hF951]=8'hF4; mem['hF952]=8'h9F; mem['hF953]=8'h83;
    mem['hF954]=8'h7E; mem['hF955]=8'hE4; mem['hF956]=8'h4B; mem['hF957]=8'h81;
    mem['hF958]=8'h45; mem['hF959]=8'h27; mem['hF95A]=8'hF1; mem['hF95B]=8'h81;
    mem['hF95C]=8'h51; mem['hF95D]=8'h26; mem['hF95E]=8'h06; mem['hF95F]=8'hBD;
    mem['hF960]=8'hF0; mem['hF961]=8'hA2; mem['hF962]=8'h7E; mem['hF963]=8'hE4;
    mem['hF964]=8'h22; mem['hF965]=8'h8D; mem['hF966]=8'h02; mem['hF967]=8'h20;
    mem['hF968]=8'hAD; mem['hF969]=8'h81; mem['hF96A]=8'h20; mem['hF96B]=8'h26;
    mem['hF96C]=8'h10; mem['hF96D]=8'h8C; mem['hF96E]=8'hC6; mem['hF96F]=8'hF9;
    mem['hF970]=8'hA6; mem['hF971]=8'h84; mem['hF972]=8'h27; mem['hF973]=8'h08;
    mem['hF974]=8'hBD; mem['hF975]=8'hE0; mem['hF976]=8'h14; mem['hF977]=8'h30;
    mem['hF978]=8'h01; mem['hF979]=8'h5A; mem['hF97A]=8'h26; mem['hF97B]=8'hF4;
    mem['hF97C]=8'h39; mem['hF97D]=8'h81; mem['hF97E]=8'h44; mem['hF97F]=8'h26;
    mem['hF980]=8'h48; mem['hF981]=8'h6D; mem['hF982]=8'h84; mem['hF983]=8'h27;
    mem['hF984]=8'hF7; mem['hF985]=8'h8D; mem['hF986]=8'h04; mem['hF987]=8'h5A;
    mem['hF988]=8'h26; mem['hF989]=8'hF7; mem['hF98A]=8'h39; mem['hF98B]=8'h0A;
    mem['hF98C]=8'h97; mem['hF98D]=8'h31; mem['hF98E]=8'h1F; mem['hF98F]=8'h31;
    mem['hF990]=8'h21; mem['hF991]=8'hA6; mem['hF992]=8'h21; mem['hF993]=8'hA7;
    mem['hF994]=8'hA4; mem['hF995]=8'h26; mem['hF996]=8'hF8; mem['hF997]=8'h39;
    mem['hF998]=8'h81; mem['hF999]=8'h49; mem['hF99A]=8'h27; mem['hF99B]=8'h13;
    mem['hF99C]=8'h81; mem['hF99D]=8'h58; mem['hF99E]=8'h27; mem['hF99F]=8'h0D;
    mem['hF9A0]=8'h81; mem['hF9A1]=8'h48; mem['hF9A2]=8'h26; mem['hF9A3]=8'h5C;
    mem['hF9A4]=8'h6F; mem['hF9A5]=8'h84; mem['hF9A6]=8'h1F; mem['hF9A7]=8'h10;
    mem['hF9A8]=8'h83; mem['hF9A9]=8'h00; mem['hF9AA]=8'hF5; mem['hF9AB]=8'hD7;
    mem['hF9AC]=8'h97; mem['hF9AD]=8'h8D; mem['hF9AE]=8'hBF; mem['hF9AF]=8'hBD;
    mem['hF9B0]=8'hFA; mem['hF9B1]=8'h41; mem['hF9B2]=8'h81; mem['hF9B3]=8'h0D;
    mem['hF9B4]=8'h27; mem['hF9B5]=8'h8E; mem['hF9B6]=8'h81; mem['hF9B7]=8'h1B;
    mem['hF9B8]=8'h27; mem['hF9B9]=8'h25; mem['hF9BA]=8'h81; mem['hF9BB]=8'h08;
    mem['hF9BC]=8'h26; mem['hF9BD]=8'h22; mem['hF9BE]=8'h8C; mem['hF9BF]=8'h00;
    mem['hF9C0]=8'hF4; mem['hF9C1]=8'h27; mem['hF9C2]=8'hEC; mem['hF9C3]=8'h8D;
    mem['hF9C4]=8'h45; mem['hF9C5]=8'h8D; mem['hF9C6]=8'hC4; mem['hF9C7]=8'h20;
    mem['hF9C8]=8'hE6; mem['hF9C9]=8'h81; mem['hF9CA]=8'h43; mem['hF9CB]=8'h26;
    mem['hF9CC]=8'hCB; mem['hF9CD]=8'h6D; mem['hF9CE]=8'h84; mem['hF9CF]=8'h27;
    mem['hF9D0]=8'h0E; mem['hF9D1]=8'hBD; mem['hF9D2]=8'hFA; mem['hF9D3]=8'h41;
    mem['hF9D4]=8'h25; mem['hF9D5]=8'h02; mem['hF9D6]=8'h20; mem['hF9D7]=8'hF5;
    mem['hF9D8]=8'hA7; mem['hF9D9]=8'h80; mem['hF9DA]=8'h8D; mem['hF9DB]=8'h37;
    mem['hF9DC]=8'h5A; mem['hF9DD]=8'h26; mem['hF9DE]=8'hEE; mem['hF9DF]=8'h39;
    mem['hF9E0]=8'hD6; mem['hF9E1]=8'h97; mem['hF9E2]=8'hC1; mem['hF9E3]=8'hF9;
    mem['hF9E4]=8'h26; mem['hF9E5]=8'h02; mem['hF9E6]=8'h20; mem['hF9E7]=8'hC7;
    mem['hF9E8]=8'h34; mem['hF9E9]=8'h10; mem['hF9EA]=8'h6D; mem['hF9EB]=8'h80;
    mem['hF9EC]=8'h26; mem['hF9ED]=8'hFC; mem['hF9EE]=8'hE6; mem['hF9EF]=8'h82;
    mem['hF9F0]=8'hE7; mem['hF9F1]=8'h01; mem['hF9F2]=8'hAC; mem['hF9F3]=8'hE4;
    mem['hF9F4]=8'h26; mem['hF9F5]=8'hF8; mem['hF9F6]=8'h32; mem['hF9F7]=8'h62;
    mem['hF9F8]=8'hA7; mem['hF9F9]=8'h80; mem['hF9FA]=8'h8D; mem['hF9FB]=8'h17;
    mem['hF9FC]=8'h0C; mem['hF9FD]=8'h97; mem['hF9FE]=8'h20; mem['hF9FF]=8'hAF;
    mem['hFA00]=8'h81; mem['hFA01]=8'h08; mem['hFA02]=8'h26; mem['hFA03]=8'h12;
    mem['hFA04]=8'h8D; mem['hFA05]=8'h04; mem['hFA06]=8'h5A; mem['hFA07]=8'h26;
    mem['hFA08]=8'hFB; mem['hFA09]=8'h39; mem['hFA0A]=8'h8C; mem['hFA0B]=8'h00;
    mem['hFA0C]=8'hF4; mem['hFA0D]=8'h27; mem['hFA0E]=8'hD0; mem['hFA0F]=8'h30;
    mem['hFA10]=8'h1F; mem['hFA11]=8'h86; mem['hFA12]=8'h08; mem['hFA13]=8'h7E;
    mem['hFA14]=8'hE0; mem['hFA15]=8'h14; mem['hFA16]=8'h81; mem['hFA17]=8'h4B;
    mem['hFA18]=8'h27; mem['hFA19]=8'h05; mem['hFA1A]=8'h80; mem['hFA1B]=8'h53;
    mem['hFA1C]=8'h27; mem['hFA1D]=8'h01; mem['hFA1E]=8'h39; mem['hFA1F]=8'h34;
    mem['hFA20]=8'h02; mem['hFA21]=8'h8D; mem['hFA22]=8'h1E; mem['hFA23]=8'h34;
    mem['hFA24]=8'h02; mem['hFA25]=8'hA6; mem['hFA26]=8'h84; mem['hFA27]=8'h27;
    mem['hFA28]=8'h16; mem['hFA29]=8'h6D; mem['hFA2A]=8'h61; mem['hFA2B]=8'h26;
    mem['hFA2C]=8'h06; mem['hFA2D]=8'h8D; mem['hFA2E]=8'hE4; mem['hFA2F]=8'h30;
    mem['hFA30]=8'h01; mem['hFA31]=8'h20; mem['hFA32]=8'h03; mem['hFA33]=8'hBD;
    mem['hFA34]=8'hF9; mem['hFA35]=8'h8B; mem['hFA36]=8'hA6; mem['hFA37]=8'h84;
    mem['hFA38]=8'hA1; mem['hFA39]=8'hE4; mem['hFA3A]=8'h26; mem['hFA3B]=8'hE9;
    mem['hFA3C]=8'h5A; mem['hFA3D]=8'h26; mem['hFA3E]=8'hE6; mem['hFA3F]=8'h35;
    mem['hFA40]=8'hA0; mem['hFA41]=8'hBD; mem['hFA42]=8'hE0; mem['hFA43]=8'h00;
    mem['hFA44]=8'h81; mem['hFA45]=8'h7F; mem['hFA46]=8'h24; mem['hFA47]=8'hF9;
    mem['hFA48]=8'h81; mem['hFA49]=8'h5F; mem['hFA4A]=8'h26; mem['hFA4B]=8'h02;
    mem['hFA4C]=8'h86; mem['hFA4D]=8'h1B; mem['hFA4E]=8'h81; mem['hFA4F]=8'h0D;
    mem['hFA50]=8'h27; mem['hFA51]=8'h0E; mem['hFA52]=8'h81; mem['hFA53]=8'h1B;
    mem['hFA54]=8'h27; mem['hFA55]=8'h0A; mem['hFA56]=8'h81; mem['hFA57]=8'h08;
    mem['hFA58]=8'h27; mem['hFA59]=8'h06; mem['hFA5A]=8'h81; mem['hFA5B]=8'h20;
    mem['hFA5C]=8'h25; mem['hFA5D]=8'hE3; mem['hFA5E]=8'h1A; mem['hFA5F]=8'h01;
    mem['hFA60]=8'h39; mem['hFA61]=8'h86; mem['hFA62]=8'h4F; mem['hFA63]=8'h97;
    mem['hFA64]=8'h8C; mem['hFA65]=8'h39; mem['hFA66]=8'h86; mem['hFA67]=8'h00;
    mem['hFA68]=8'hD6; mem['hFA69]=8'h79; mem['hFA6A]=8'h1D; mem['hFA6B]=8'h7E;
    mem['hFA6C]=8'hEC; mem['hFA6D]=8'h78; mem['hFA6E]=8'hBD; mem['hFA6F]=8'hE9;
    mem['hFA70]=8'hF3; mem['hFA71]=8'hDC; mem['hFA72]=8'h1F; mem['hFA73]=8'h34;
    mem['hFA74]=8'h06; mem['hFA75]=8'hBD; mem['hFA76]=8'hEA; mem['hFA77]=8'hDB;
    mem['hFA78]=8'hBD; mem['hFA79]=8'hE9; mem['hFA7A]=8'hF0; mem['hFA7B]=8'h35;
    mem['hFA7C]=8'h06; mem['hFA7D]=8'h1E; mem['hFA7E]=8'h10; mem['hFA7F]=8'h9C;
    mem['hFA80]=8'h1F; mem['hFA81]=8'h26; mem['hFA82]=8'h51; mem['hFA83]=8'h7E;
    mem['hFA84]=8'hEC; mem['hFA85]=8'h78; mem['hFA86]=8'h9D; mem['hFA87]=8'h7C;
    mem['hFA88]=8'hBD; mem['hFA89]=8'hE9; mem['hFA8A]=8'hF3; mem['hFA8B]=8'hBD;
    mem['hFA8C]=8'hEA; mem['hFA8D]=8'hDB; mem['hFA8E]=8'h34; mem['hFA8F]=8'h10;
    mem['hFA90]=8'hEC; mem['hFA91]=8'h02; mem['hFA92]=8'h10; mem['hFA93]=8'h93;
    mem['hFA94]=8'h21; mem['hFA95]=8'h23; mem['hFA96]=8'h04; mem['hFA97]=8'h93;
    mem['hFA98]=8'h27; mem['hFA99]=8'h23; mem['hFA9A]=8'h12; mem['hFA9B]=8'hE6;
    mem['hFA9C]=8'h84; mem['hFA9D]=8'hBD; mem['hFA9E]=8'hEC; mem['hFA9F]=8'hF1;
    mem['hFAA0]=8'h34; mem['hFAA1]=8'h10; mem['hFAA2]=8'hAE; mem['hFAA3]=8'h62;
    mem['hFAA4]=8'hBD; mem['hFAA5]=8'hED; mem['hFAA6]=8'hC7; mem['hFAA7]=8'h35;
    mem['hFAA8]=8'h50; mem['hFAA9]=8'hAF; mem['hFAAA]=8'h42; mem['hFAAB]=8'h34;
    mem['hFAAC]=8'h40; mem['hFAAD]=8'hBD; mem['hFAAE]=8'hEE; mem['hFAAF]=8'hBC;
    mem['hFAB0]=8'h34; mem['hFAB1]=8'h04; mem['hFAB2]=8'h5D; mem['hFAB3]=8'h27;
    mem['hFAB4]=8'h1F; mem['hFAB5]=8'hC6; mem['hFAB6]=8'hFF; mem['hFAB7]=8'h81;
    mem['hFAB8]=8'h29; mem['hFAB9]=8'h27; mem['hFABA]=8'h03; mem['hFABB]=8'hBD;
    mem['hFABC]=8'hEE; mem['hFABD]=8'hBC; mem['hFABE]=8'h34; mem['hFABF]=8'h04;
    mem['hFAC0]=8'hBD; mem['hFAC1]=8'hE9; mem['hFAC2]=8'hF0; mem['hFAC3]=8'hC6;
    mem['hFAC4]=8'hAE; mem['hFAC5]=8'hBD; mem['hFAC6]=8'hE9; mem['hFAC7]=8'hF8;
    mem['hFAC8]=8'h8D; mem['hFAC9]=8'h2E; mem['hFACA]=8'h1F; mem['hFACB]=8'h13;
    mem['hFACC]=8'hAE; mem['hFACD]=8'h62; mem['hFACE]=8'hA6; mem['hFACF]=8'h84;
    mem['hFAD0]=8'hA0; mem['hFAD1]=8'h61; mem['hFAD2]=8'h24; mem['hFAD3]=8'h03;
    mem['hFAD4]=8'h7E; mem['hFAD5]=8'hEB; mem['hFAD6]=8'hCE; mem['hFAD7]=8'h4C;
    mem['hFAD8]=8'hA1; mem['hFAD9]=8'hE4; mem['hFADA]=8'h24; mem['hFADB]=8'h02;
    mem['hFADC]=8'hA7; mem['hFADD]=8'hE4; mem['hFADE]=8'hA6; mem['hFADF]=8'h61;
    mem['hFAE0]=8'h1E; mem['hFAE1]=8'h89; mem['hFAE2]=8'hAE; mem['hFAE3]=8'h02;
    mem['hFAE4]=8'h5A; mem['hFAE5]=8'h3A; mem['hFAE6]=8'h4D; mem['hFAE7]=8'h27;
    mem['hFAE8]=8'h0D; mem['hFAE9]=8'hA1; mem['hFAEA]=8'hE4; mem['hFAEB]=8'h23;
    mem['hFAEC]=8'h02; mem['hFAED]=8'hA6; mem['hFAEE]=8'hE4; mem['hFAEF]=8'h1F;
    mem['hFAF0]=8'h89; mem['hFAF1]=8'h1E; mem['hFAF2]=8'h31; mem['hFAF3]=8'hBD;
    mem['hFAF4]=8'hE1; mem['hFAF5]=8'hAE; mem['hFAF6]=8'h35; mem['hFAF7]=8'h96;
    mem['hFAF8]=8'hBD; mem['hFAF9]=8'hE8; mem['hFAFA]=8'hDF; mem['hFAFB]=8'h7E;
    mem['hFAFC]=8'hED; mem['hFAFD]=8'hD8; mem['hFAFE]=8'hBD; mem['hFAFF]=8'hE9;
    mem['hFB00]=8'hF3; mem['hFB01]=8'hBD; mem['hFB02]=8'hEE; mem['hFB03]=8'h8F;
    mem['hFB04]=8'h34; mem['hFB05]=8'h04; mem['hFB06]=8'hBD; mem['hFB07]=8'hE9;
    mem['hFB08]=8'hF6; mem['hFB09]=8'hBD; mem['hFB0A]=8'hE8; mem['hFB0B]=8'hDF;
    mem['hFB0C]=8'hBD; mem['hFB0D]=8'hE9; mem['hFB0E]=8'hF0; mem['hFB0F]=8'h96;
    mem['hFB10]=8'h06; mem['hFB11]=8'h26; mem['hFB12]=8'h05; mem['hFB13]=8'hBD;
    mem['hFB14]=8'hEE; mem['hFB15]=8'h92; mem['hFB16]=8'h20; mem['hFB17]=8'h03;
    mem['hFB18]=8'hBD; mem['hFB19]=8'hEE; mem['hFB1A]=8'h28; mem['hFB1B]=8'h34;
    mem['hFB1C]=8'h04; mem['hFB1D]=8'hE6; mem['hFB1E]=8'h61; mem['hFB1F]=8'hBD;
    mem['hFB20]=8'hEC; mem['hFB21]=8'h93; mem['hFB22]=8'h35; mem['hFB23]=8'h06;
    mem['hFB24]=8'h27; mem['hFB25]=8'h05; mem['hFB26]=8'hA7; mem['hFB27]=8'h80;
    mem['hFB28]=8'h5A; mem['hFB29]=8'h26; mem['hFB2A]=8'hFB; mem['hFB2B]=8'h7E;
    mem['hFB2C]=8'hEE; mem['hFB2D]=8'h1F; mem['hFB2E]=8'hBD; mem['hFB2F]=8'hE9;
    mem['hFB30]=8'hF3; mem['hFB31]=8'hBD; mem['hFB32]=8'hE8; mem['hFB33]=8'hDF;
    mem['hFB34]=8'hC6; mem['hFB35]=8'h01; mem['hFB36]=8'h34; mem['hFB37]=8'h04;
    mem['hFB38]=8'h96; mem['hFB39]=8'h06; mem['hFB3A]=8'h26; mem['hFB3B]=8'h10;
    mem['hFB3C]=8'hBD; mem['hFB3D]=8'hEE; mem['hFB3E]=8'h92; mem['hFB3F]=8'hE7;
    mem['hFB40]=8'hE4; mem['hFB41]=8'h27; mem['hFB42]=8'h91; mem['hFB43]=8'hBD;
    mem['hFB44]=8'hE9; mem['hFB45]=8'hF6; mem['hFB46]=8'hBD; mem['hFB47]=8'hE8;
    mem['hFB48]=8'hDF; mem['hFB49]=8'hBD; mem['hFB4A]=8'hE8; mem['hFB4B]=8'hCF;
    mem['hFB4C]=8'h9E; mem['hFB4D]=8'h52; mem['hFB4E]=8'h34; mem['hFB4F]=8'h10;
    mem['hFB50]=8'hBD; mem['hFB51]=8'hE9; mem['hFB52]=8'hF6; mem['hFB53]=8'hBD;
    mem['hFB54]=8'hFA; mem['hFB55]=8'hF8; mem['hFB56]=8'h34; mem['hFB57]=8'h14;
    mem['hFB58]=8'hBD; mem['hFB59]=8'hE9; mem['hFB5A]=8'hF0; mem['hFB5B]=8'hAE;
    mem['hFB5C]=8'h63; mem['hFB5D]=8'hBD; mem['hFB5E]=8'hED; mem['hFB5F]=8'hDD;
    mem['hFB60]=8'h34; mem['hFB61]=8'h04; mem['hFB62]=8'hE1; mem['hFB63]=8'h66;
    mem['hFB64]=8'h25; mem['hFB65]=8'h23; mem['hFB66]=8'hA6; mem['hFB67]=8'h61;
    mem['hFB68]=8'h27; mem['hFB69]=8'h1C; mem['hFB6A]=8'hE6; mem['hFB6B]=8'h66;
    mem['hFB6C]=8'h5A; mem['hFB6D]=8'h3A; mem['hFB6E]=8'h31; mem['hFB6F]=8'h84;
    mem['hFB70]=8'hEE; mem['hFB71]=8'h62; mem['hFB72]=8'hE6; mem['hFB73]=8'h61;
    mem['hFB74]=8'hA6; mem['hFB75]=8'hE4; mem['hFB76]=8'hA0; mem['hFB77]=8'h66;
    mem['hFB78]=8'h4C; mem['hFB79]=8'hA1; mem['hFB7A]=8'h61; mem['hFB7B]=8'h25;
    mem['hFB7C]=8'h0C; mem['hFB7D]=8'hA6; mem['hFB7E]=8'h80; mem['hFB7F]=8'hA1;
    mem['hFB80]=8'hC0; mem['hFB81]=8'h26; mem['hFB82]=8'h0C; mem['hFB83]=8'h5A;
    mem['hFB84]=8'h26; mem['hFB85]=8'hF7; mem['hFB86]=8'hE6; mem['hFB87]=8'h66;
    mem['hFB88]=8'h21; mem['hFB89]=8'h5F; mem['hFB8A]=8'h32; mem['hFB8B]=8'h67;
    mem['hFB8C]=8'h7E; mem['hFB8D]=8'hEC; mem['hFB8E]=8'h77; mem['hFB8F]=8'h6C;
    mem['hFB90]=8'h66; mem['hFB91]=8'h30; mem['hFB92]=8'h21; mem['hFB93]=8'h20;
    mem['hFB94]=8'hD9; mem['hFB95]=8'h81; mem['hFB96]=8'h26; mem['hFB97]=8'h26;
    mem['hFB98]=8'h5C; mem['hFB99]=8'h32; mem['hFB9A]=8'h62; mem['hFB9B]=8'h0F;
    mem['hFB9C]=8'h52; mem['hFB9D]=8'h0F; mem['hFB9E]=8'h53; mem['hFB9F]=8'h8E;
    mem['hFBA0]=8'h00; mem['hFBA1]=8'h52; mem['hFBA2]=8'h9D; mem['hFBA3]=8'h7C;
    mem['hFBA4]=8'h81; mem['hFBA5]=8'h4F; mem['hFBA6]=8'h27; mem['hFBA7]=8'h12;
    mem['hFBA8]=8'h81; mem['hFBA9]=8'h48; mem['hFBAA]=8'h27; mem['hFBAB]=8'h23;
    mem['hFBAC]=8'h9D; mem['hFBAD]=8'h82; mem['hFBAE]=8'h20; mem['hFBAF]=8'h0C;
    mem['hFBB0]=8'h81; mem['hFBB1]=8'h38; mem['hFBB2]=8'h10; mem['hFBB3]=8'h22;
    mem['hFBB4]=8'hEE; mem['hFBB5]=8'h4A; mem['hFBB6]=8'hC6; mem['hFBB7]=8'h03;
    mem['hFBB8]=8'h8D; mem['hFBB9]=8'h2A; mem['hFBBA]=8'h9D; mem['hFBBB]=8'h7C;
    mem['hFBBC]=8'h25; mem['hFBBD]=8'hF2; mem['hFBBE]=8'h0F; mem['hFBBF]=8'h50;
    mem['hFBC0]=8'h0F; mem['hFBC1]=8'h51; mem['hFBC2]=8'h0F; mem['hFBC3]=8'h06;
    mem['hFBC4]=8'h0F; mem['hFBC5]=8'h63; mem['hFBC6]=8'h0F; mem['hFBC7]=8'h54;
    mem['hFBC8]=8'hC6; mem['hFBC9]=8'hA0; mem['hFBCA]=8'hD7; mem['hFBCB]=8'h4F;
    mem['hFBCC]=8'h7E; mem['hFBCD]=8'hF1; mem['hFBCE]=8'h62; mem['hFBCF]=8'h9D;
    mem['hFBD0]=8'h7C; mem['hFBD1]=8'h25; mem['hFBD2]=8'h0B; mem['hFBD3]=8'hBD;
    mem['hFBD4]=8'hEB; mem['hFBD5]=8'h26; mem['hFBD6]=8'h25; mem['hFBD7]=8'hE6;
    mem['hFBD8]=8'h81; mem['hFBD9]=8'h47; mem['hFBDA]=8'h24; mem['hFBDB]=8'hE2;
    mem['hFBDC]=8'h80; mem['hFBDD]=8'h07; mem['hFBDE]=8'hC6; mem['hFBDF]=8'h04;
    mem['hFBE0]=8'h8D; mem['hFBE1]=8'h02; mem['hFBE2]=8'h20; mem['hFBE3]=8'hEB;
    mem['hFBE4]=8'h68; mem['hFBE5]=8'h01; mem['hFBE6]=8'h69; mem['hFBE7]=8'h84;
    mem['hFBE8]=8'h10; mem['hFBE9]=8'h25; mem['hFBEA]=8'hF5; mem['hFBEB]=8'hEC;
    mem['hFBEC]=8'h5A; mem['hFBED]=8'h26; mem['hFBEE]=8'hF5; mem['hFBEF]=8'h80;
    mem['hFBF0]=8'h30; mem['hFBF1]=8'hAB; mem['hFBF2]=8'h01; mem['hFBF3]=8'hA7;
    mem['hFBF4]=8'h01; mem['hFBF5]=8'h39; mem['hFBF6]=8'h35; mem['hFBF7]=8'h40;
    mem['hFBF8]=8'h0F; mem['hFBF9]=8'h06; mem['hFBFA]=8'h9E; mem['hFBFB]=8'h83;
    mem['hFBFC]=8'h9D; mem['hFBFD]=8'h7C; mem['hFBFE]=8'h81; mem['hFBFF]=8'h26;
    mem['hFC00]=8'h27; mem['hFC01]=8'h99; mem['hFC02]=8'h81; mem['hFC03]=8'hB0;
    mem['hFC04]=8'h27; mem['hFC05]=8'h5E; mem['hFC06]=8'h81; mem['hFC07]=8'hFF;
    mem['hFC08]=8'h26; mem['hFC09]=8'h08; mem['hFC0A]=8'h9D; mem['hFC0B]=8'h7C;
    mem['hFC0C]=8'h81; mem['hFC0D]=8'h83; mem['hFC0E]=8'h10; mem['hFC0F]=8'h27;
    mem['hFC10]=8'h00; mem['hFC11]=8'hAB; mem['hFC12]=8'h9F; mem['hFC13]=8'h83;
    mem['hFC14]=8'h6E; mem['hFC15]=8'hC4; mem['hFC16]=8'h9E; mem['hFC17]=8'h68;
    mem['hFC18]=8'h30; mem['hFC19]=8'h01; mem['hFC1A]=8'h26; mem['hFC1B]=8'hD9;
    mem['hFC1C]=8'hC6; mem['hFC1D]=8'h16; mem['hFC1E]=8'h7E; mem['hFC1F]=8'hE4;
    mem['hFC20]=8'h03; mem['hFC21]=8'hAE; mem['hFC22]=8'h9F; mem['hFC23]=8'h00;
    mem['hFC24]=8'h83; mem['hFC25]=8'h8C; mem['hFC26]=8'hFF; mem['hFC27]=8'h83;
    mem['hFC28]=8'h10; mem['hFC29]=8'h27; mem['hFC2A]=8'h00; mem['hFC2B]=8'h74;
    mem['hFC2C]=8'h8D; mem['hFC2D]=8'h23; mem['hFC2E]=8'h8D; mem['hFC2F]=8'hE6;
    mem['hFC30]=8'hBD; mem['hFC31]=8'hE9; mem['hFC32]=8'hF3; mem['hFC33]=8'hC6;
    mem['hFC34]=8'h80; mem['hFC35]=8'hD7; mem['hFC36]=8'h08; mem['hFC37]=8'hBD;
    mem['hFC38]=8'hEA; mem['hFC39]=8'hDB; mem['hFC3A]=8'h8D; mem['hFC3B]=8'h25;
    mem['hFC3C]=8'hBD; mem['hFC3D]=8'hE9; mem['hFC3E]=8'hF0; mem['hFC3F]=8'hC6;
    mem['hFC40]=8'hAE; mem['hFC41]=8'hBD; mem['hFC42]=8'hE9; mem['hFC43]=8'hF8;
    mem['hFC44]=8'h9E; mem['hFC45]=8'h4B; mem['hFC46]=8'hDC; mem['hFC47]=8'h83;
    mem['hFC48]=8'hED; mem['hFC49]=8'h84; mem['hFC4A]=8'hDC; mem['hFC4B]=8'h39;
    mem['hFC4C]=8'hED; mem['hFC4D]=8'h02; mem['hFC4E]=8'h7E; mem['hFC4F]=8'hE6;
    mem['hFC50]=8'h8D; mem['hFC51]=8'hC6; mem['hFC52]=8'hB0; mem['hFC53]=8'hBD;
    mem['hFC54]=8'hE9; mem['hFC55]=8'hF8; mem['hFC56]=8'hC6; mem['hFC57]=8'h80;
    mem['hFC58]=8'hD7; mem['hFC59]=8'h08; mem['hFC5A]=8'h8A; mem['hFC5B]=8'h80;
    mem['hFC5C]=8'hBD; mem['hFC5D]=8'hEA; mem['hFC5E]=8'hE0; mem['hFC5F]=8'h9F;
    mem['hFC60]=8'h4B; mem['hFC61]=8'h7E; mem['hFC62]=8'hE8; mem['hFC63]=8'hCC;
    mem['hFC64]=8'h8D; mem['hFC65]=8'hEB; mem['hFC66]=8'h34; mem['hFC67]=8'h10;
    mem['hFC68]=8'hBD; mem['hFC69]=8'hE9; mem['hFC6A]=8'hEB; mem['hFC6B]=8'h8D;
    mem['hFC6C]=8'hF4; mem['hFC6D]=8'h35; mem['hFC6E]=8'h40; mem['hFC6F]=8'hC6;
    mem['hFC70]=8'h32; mem['hFC71]=8'hAE; mem['hFC72]=8'h42; mem['hFC73]=8'h27;
    mem['hFC74]=8'hA9; mem['hFC75]=8'h10; mem['hFC76]=8'h9E; mem['hFC77]=8'h83;
    mem['hFC78]=8'hEE; mem['hFC79]=8'hC4; mem['hFC7A]=8'hDF; mem['hFC7B]=8'h83;
    mem['hFC7C]=8'hA6; mem['hFC7D]=8'h04; mem['hFC7E]=8'h34; mem['hFC7F]=8'h02;
    mem['hFC80]=8'hEC; mem['hFC81]=8'h84; mem['hFC82]=8'hEE; mem['hFC83]=8'h02;
    mem['hFC84]=8'h34; mem['hFC85]=8'h76; mem['hFC86]=8'hBD; mem['hFC87]=8'hF3;
    mem['hFC88]=8'h7B; mem['hFC89]=8'hBD; mem['hFC8A]=8'hE8; mem['hFC8B]=8'hCA;
    mem['hFC8C]=8'h35; mem['hFC8D]=8'h76; mem['hFC8E]=8'hED; mem['hFC8F]=8'h84;
    mem['hFC90]=8'hEF; mem['hFC91]=8'h02; mem['hFC92]=8'h35; mem['hFC93]=8'h02;
    mem['hFC94]=8'hA7; mem['hFC95]=8'h04; mem['hFC96]=8'h9D; mem['hFC97]=8'h82;
    mem['hFC98]=8'h10; mem['hFC99]=8'h26; mem['hFC9A]=8'hED; mem['hFC9B]=8'h64;
    mem['hFC9C]=8'h10; mem['hFC9D]=8'h9F; mem['hFC9E]=8'h83; mem['hFC9F]=8'h39;
    mem['hFCA0]=8'h9D; mem['hFCA1]=8'h7C; mem['hFCA2]=8'h8D; mem['hFCA3]=8'h09;
    mem['hFCA4]=8'h34; mem['hFCA5]=8'h10; mem['hFCA6]=8'h8D; mem['hFCA7]=8'h2D;
    mem['hFCA8]=8'h35; mem['hFCA9]=8'h40; mem['hFCAA]=8'hAF; mem['hFCAB]=8'hC4;
    mem['hFCAC]=8'h39; mem['hFCAD]=8'h5F; mem['hFCAE]=8'h9D; mem['hFCAF]=8'h7C;
    mem['hFCB0]=8'h24; mem['hFCB1]=8'h06; mem['hFCB2]=8'h80; mem['hFCB3]=8'h30;
    mem['hFCB4]=8'h1F; mem['hFCB5]=8'h89; mem['hFCB6]=8'h9D; mem['hFCB7]=8'h7C;
    mem['hFCB8]=8'h9E; mem['hFCB9]=8'h8D; mem['hFCBA]=8'h58; mem['hFCBB]=8'h3A;
    mem['hFCBC]=8'h39; mem['hFCBD]=8'h8D; mem['hFCBE]=8'hEE; mem['hFCBF]=8'hAE;
    mem['hFCC0]=8'h84; mem['hFCC1]=8'h34; mem['hFCC2]=8'h10; mem['hFCC3]=8'hBD;
    mem['hFCC4]=8'hE9; mem['hFCC5]=8'hEB; mem['hFCC6]=8'h8E; mem['hFCC7]=8'h00;
    mem['hFCC8]=8'h4F; mem['hFCC9]=8'h96; mem['hFCCA]=8'h06; mem['hFCCB]=8'h27;
    mem['hFCCC]=8'h07; mem['hFCCD]=8'hBD; mem['hFCCE]=8'hED; mem['hFCCF]=8'hDB;
    mem['hFCD0]=8'h9E; mem['hFCD1]=8'h52; mem['hFCD2]=8'h96; mem['hFCD3]=8'h06;
    mem['hFCD4]=8'h39; mem['hFCD5]=8'hC6; mem['hFCD6]=8'hAE; mem['hFCD7]=8'hBD;
    mem['hFCD8]=8'hE9; mem['hFCD9]=8'hF8; mem['hFCDA]=8'h7E; mem['hFCDB]=8'hEE;
    mem['hFCDC]=8'hC1; mem['hFCDD]=8'h10; mem['hFCDE]=8'h27; mem['hFCDF]=8'hEE;
    mem['hFCE0]=8'hED; mem['hFCE1]=8'hBD; mem['hFCE2]=8'hE7; mem['hFCE3]=8'h14;
    mem['hFCE4]=8'hBD; mem['hFCE5]=8'hE4; mem['hFCE6]=8'hA2; mem['hFCE7]=8'h9F;
    mem['hFCE8]=8'h93; mem['hFCE9]=8'h9D; mem['hFCEA]=8'h82; mem['hFCEB]=8'h27;
    mem['hFCEC]=8'h10; mem['hFCED]=8'h81; mem['hFCEE]=8'hA7; mem['hFCEF]=8'h26;
    mem['hFCF0]=8'h3B; mem['hFCF1]=8'h9D; mem['hFCF2]=8'h7C; mem['hFCF3]=8'h27;
    mem['hFCF4]=8'h04; mem['hFCF5]=8'h8D; mem['hFCF6]=8'h24; mem['hFCF7]=8'h20;
    mem['hFCF8]=8'h04; mem['hFCF9]=8'h86; mem['hFCFA]=8'hFF; mem['hFCFB]=8'h97;
    mem['hFCFC]=8'h2B; mem['hFCFD]=8'hDE; mem['hFCFE]=8'h93; mem['hFCFF]=8'h8C;
    mem['hFD00]=8'hEE; mem['hFD01]=8'hC4; mem['hFD02]=8'hEC; mem['hFD03]=8'hC4;
    mem['hFD04]=8'h27; mem['hFD05]=8'h06; mem['hFD06]=8'hEC; mem['hFD07]=8'h42;
    mem['hFD08]=8'h93; mem['hFD09]=8'h2B; mem['hFD0A]=8'h23; mem['hFD0B]=8'hF4;
    mem['hFD0C]=8'h9E; mem['hFD0D]=8'h93; mem['hFD0E]=8'h8D; mem['hFD0F]=8'h15;
    mem['hFD10]=8'hBD; mem['hFD11]=8'hE4; mem['hFD12]=8'hC2; mem['hFD13]=8'h9E;
    mem['hFD14]=8'h93; mem['hFD15]=8'hBD; mem['hFD16]=8'hE4; mem['hFD17]=8'h92;
    mem['hFD18]=8'h7E; mem['hFD19]=8'hE4; mem['hFD1A]=8'h22; mem['hFD1B]=8'hBD;
    mem['hFD1C]=8'hE7; mem['hFD1D]=8'h14; mem['hFD1E]=8'h7E; mem['hFD1F]=8'hE1;
    mem['hFD20]=8'hB7; mem['hFD21]=8'hA6; mem['hFD22]=8'hC0; mem['hFD23]=8'hA7;
    mem['hFD24]=8'h80; mem['hFD25]=8'h11; mem['hFD26]=8'h93; mem['hFD27]=8'h1B;
    mem['hFD28]=8'h26; mem['hFD29]=8'hF7; mem['hFD2A]=8'h9F; mem['hFD2B]=8'h1B;
    mem['hFD2C]=8'h39; mem['hFD2D]=8'hBD; mem['hFD2E]=8'hFC; mem['hFD2F]=8'h16;
    mem['hFD30]=8'h9D; mem['hFD31]=8'h7C; mem['hFD32]=8'h81; mem['hFD33]=8'h22;
    mem['hFD34]=8'h26; mem['hFD35]=8'h0B; mem['hFD36]=8'hBD; mem['hFD37]=8'hE9;
    mem['hFD38]=8'hCD; mem['hFD39]=8'hC6; mem['hFD3A]=8'h3B; mem['hFD3B]=8'hBD;
    mem['hFD3C]=8'hE9; mem['hFD3D]=8'hF8; mem['hFD3E]=8'hBD; mem['hFD3F]=8'hF0;
    mem['hFD40]=8'hE5; mem['hFD41]=8'h32; mem['hFD42]=8'h7E; mem['hFD43]=8'hBD;
    mem['hFD44]=8'hE7; mem['hFD45]=8'hC9; mem['hFD46]=8'h32; mem['hFD47]=8'h62;
    mem['hFD48]=8'hBD; mem['hFD49]=8'hEA; mem['hFD4A]=8'hDB; mem['hFD4B]=8'h9F;
    mem['hFD4C]=8'h3B; mem['hFD4D]=8'hBD; mem['hFD4E]=8'hE8; mem['hFD4F]=8'hCF;
    mem['hFD50]=8'h8E; mem['hFD51]=8'h00; mem['hFD52]=8'hF3; mem['hFD53]=8'h4F;
    mem['hFD54]=8'hBD; mem['hFD55]=8'hEC; mem['hFD56]=8'hA0; mem['hFD57]=8'h7E;
    mem['hFD58]=8'hE7; mem['hFD59]=8'h51; mem['hFD5A]=8'hBD; mem['hFD5B]=8'hE7;
    mem['hFD5C]=8'h14; mem['hFD5D]=8'h9E; mem['hFD5E]=8'h2B; mem['hFD5F]=8'h39;
    mem['hFD60]=8'h9E; mem['hFD61]=8'h91; mem['hFD62]=8'h9F; mem['hFD63]=8'h2B;
    mem['hFD64]=8'h7E; mem['hFD65]=8'hE4; mem['hFD66]=8'hA2; mem['hFD67]=8'hBD;
    mem['hFD68]=8'hE4; mem['hFD69]=8'hC7; mem['hFD6A]=8'hCC; mem['hFD6B]=8'h00;
    mem['hFD6C]=8'h0A; mem['hFD6D]=8'hDD; mem['hFD6E]=8'h95; mem['hFD6F]=8'hDD;
    mem['hFD70]=8'h8F; mem['hFD71]=8'h5F; mem['hFD72]=8'hDD; mem['hFD73]=8'h91;
    mem['hFD74]=8'h9D; mem['hFD75]=8'h82; mem['hFD76]=8'h24; mem['hFD77]=8'h06;
    mem['hFD78]=8'h8D; mem['hFD79]=8'hE0; mem['hFD7A]=8'h9F; mem['hFD7B]=8'h95;
    mem['hFD7C]=8'h9D; mem['hFD7D]=8'h82; mem['hFD7E]=8'h27; mem['hFD7F]=8'h1B;
    mem['hFD80]=8'hBD; mem['hFD81]=8'hE9; mem['hFD82]=8'hF6; mem['hFD83]=8'h24;
    mem['hFD84]=8'h06; mem['hFD85]=8'h8D; mem['hFD86]=8'hD3; mem['hFD87]=8'h9F;
    mem['hFD88]=8'h91; mem['hFD89]=8'h9D; mem['hFD8A]=8'h82; mem['hFD8B]=8'h27;
    mem['hFD8C]=8'h0E; mem['hFD8D]=8'hBD; mem['hFD8E]=8'hE9; mem['hFD8F]=8'hF6;
    mem['hFD90]=8'h24; mem['hFD91]=8'h06; mem['hFD92]=8'h8D; mem['hFD93]=8'hC6;
    mem['hFD94]=8'h9F; mem['hFD95]=8'h8F; mem['hFD96]=8'h27; mem['hFD97]=8'h49;
    mem['hFD98]=8'hBD; mem['hFD99]=8'hE1; mem['hFD9A]=8'hB7; mem['hFD9B]=8'h8D;
    mem['hFD9C]=8'hC3; mem['hFD9D]=8'h9F; mem['hFD9E]=8'h93; mem['hFD9F]=8'h9E;
    mem['hFDA0]=8'h95; mem['hFDA1]=8'h8D; mem['hFDA2]=8'hBF; mem['hFDA3]=8'h9C;
    mem['hFDA4]=8'h93; mem['hFDA5]=8'h25; mem['hFDA6]=8'h3A; mem['hFDA7]=8'h8D;
    mem['hFDA8]=8'h1C; mem['hFDA9]=8'hBD; mem['hFDAA]=8'hFE; mem['hFDAB]=8'h3B;
    mem['hFDAC]=8'hBD; mem['hFDAD]=8'hE4; mem['hFDAE]=8'h90; mem['hFDAF]=8'h8D;
    mem['hFDB0]=8'hAF; mem['hFDB1]=8'h9F; mem['hFDB2]=8'h93; mem['hFDB3]=8'h8D;
    mem['hFDB4]=8'h3A; mem['hFDB5]=8'h8D; mem['hFDB6]=8'h0F; mem['hFDB7]=8'h8D;
    mem['hFDB8]=8'h36; mem['hFDB9]=8'hBD; mem['hFDBA]=8'hFE; mem['hFDBB]=8'hD6;
    mem['hFDBC]=8'hBD; mem['hFDBD]=8'hE4; mem['hFDBE]=8'hC7; mem['hFDBF]=8'hBD;
    mem['hFDC0]=8'hE4; mem['hFDC1]=8'h90; mem['hFDC2]=8'h7E; mem['hFDC3]=8'hE4;
    mem['hFDC4]=8'h22; mem['hFDC5]=8'h86; mem['hFDC6]=8'h4F; mem['hFDC7]=8'h97;
    mem['hFDC8]=8'h98; mem['hFDC9]=8'h9E; mem['hFDCA]=8'h93; mem['hFDCB]=8'hDC;
    mem['hFDCC]=8'h95; mem['hFDCD]=8'h8D; mem['hFDCE]=8'h15; mem['hFDCF]=8'h0D;
    mem['hFDD0]=8'h98; mem['hFDD1]=8'h26; mem['hFDD2]=8'h02; mem['hFDD3]=8'hED;
    mem['hFDD4]=8'h02; mem['hFDD5]=8'hAE; mem['hFDD6]=8'h84; mem['hFDD7]=8'h8D;
    mem['hFDD8]=8'h0B; mem['hFDD9]=8'hD3; mem['hFDDA]=8'h8F; mem['hFDDB]=8'h25;
    mem['hFDDC]=8'h04; mem['hFDDD]=8'h81; mem['hFDDE]=8'hFA; mem['hFDDF]=8'h25;
    mem['hFDE0]=8'hEE; mem['hFDE1]=8'h7E; mem['hFDE2]=8'hEB; mem['hFDE3]=8'hCE;
    mem['hFDE4]=8'h34; mem['hFDE5]=8'h06; mem['hFDE6]=8'hEC; mem['hFDE7]=8'h84;
    mem['hFDE8]=8'h35; mem['hFDE9]=8'h06; mem['hFDEA]=8'h26; mem['hFDEB]=8'h02;
    mem['hFDEC]=8'h32; mem['hFDED]=8'h62; mem['hFDEE]=8'h39; mem['hFDEF]=8'h9E;
    mem['hFDF0]=8'h19; mem['hFDF1]=8'h30; mem['hFDF2]=8'h1F; mem['hFDF3]=8'h30;
    mem['hFDF4]=8'h01; mem['hFDF5]=8'h8D; mem['hFDF6]=8'hED; mem['hFDF7]=8'h30;
    mem['hFDF8]=8'h03; mem['hFDF9]=8'h30; mem['hFDFA]=8'h01; mem['hFDFB]=8'hA6;
    mem['hFDFC]=8'h84; mem['hFDFD]=8'h27; mem['hFDFE]=8'hF4; mem['hFDFF]=8'h9F;
    mem['hFE00]=8'h0F; mem['hFE01]=8'h4A; mem['hFE02]=8'h27; mem['hFE03]=8'h0C;
    mem['hFE04]=8'h4A; mem['hFE05]=8'h27; mem['hFE06]=8'h2A; mem['hFE07]=8'h4A;
    mem['hFE08]=8'h26; mem['hFE09]=8'hEF; mem['hFE0A]=8'h86; mem['hFE0B]=8'h03;
    mem['hFE0C]=8'hA7; mem['hFE0D]=8'h80; mem['hFE0E]=8'h20; mem['hFE0F]=8'hE7;
    mem['hFE10]=8'hEC; mem['hFE11]=8'h01; mem['hFE12]=8'h6A; mem['hFE13]=8'h02;
    mem['hFE14]=8'h27; mem['hFE15]=8'h01; mem['hFE16]=8'h4F; mem['hFE17]=8'hE6;
    mem['hFE18]=8'h03; mem['hFE19]=8'h6A; mem['hFE1A]=8'h04; mem['hFE1B]=8'h27;
    mem['hFE1C]=8'h01; mem['hFE1D]=8'h5F; mem['hFE1E]=8'hED; mem['hFE1F]=8'h01;
    mem['hFE20]=8'hDD; mem['hFE21]=8'h2B; mem['hFE22]=8'hBD; mem['hFE23]=8'hE4;
    mem['hFE24]=8'hA2; mem['hFE25]=8'h9E; mem['hFE26]=8'h0F; mem['hFE27]=8'h25;
    mem['hFE28]=8'hE1; mem['hFE29]=8'hDC; mem['hFE2A]=8'h47; mem['hFE2B]=8'h6C;
    mem['hFE2C]=8'h80; mem['hFE2D]=8'hED; mem['hFE2E]=8'h84; mem['hFE2F]=8'h20;
    mem['hFE30]=8'hC6; mem['hFE31]=8'h6F; mem['hFE32]=8'h84; mem['hFE33]=8'hAE;
    mem['hFE34]=8'h01; mem['hFE35]=8'hAE; mem['hFE36]=8'h02; mem['hFE37]=8'h9F;
    mem['hFE38]=8'h47; mem['hFE39]=8'h20; mem['hFE3A]=8'hEA; mem['hFE3B]=8'h9E;
    mem['hFE3C]=8'h19; mem['hFE3D]=8'h20; mem['hFE3E]=8'h04; mem['hFE3F]=8'h9E;
    mem['hFE40]=8'h83; mem['hFE41]=8'h30; mem['hFE42]=8'h01; mem['hFE43]=8'h8D;
    mem['hFE44]=8'h9F; mem['hFE45]=8'h30; mem['hFE46]=8'h02; mem['hFE47]=8'h30;
    mem['hFE48]=8'h01; mem['hFE49]=8'h9F; mem['hFE4A]=8'h83; mem['hFE4B]=8'h9D;
    mem['hFE4C]=8'h7C; mem['hFE4D]=8'h4D; mem['hFE4E]=8'h27; mem['hFE4F]=8'hEF;
    mem['hFE50]=8'h2A; mem['hFE51]=8'hF9; mem['hFE52]=8'h9E; mem['hFE53]=8'h83;
    mem['hFE54]=8'h81; mem['hFE55]=8'hFF; mem['hFE56]=8'h27; mem['hFE57]=8'hEF;
    mem['hFE58]=8'h81; mem['hFE59]=8'hA2; mem['hFE5A]=8'h27; mem['hFE5B]=8'h12;
    mem['hFE5C]=8'h81; mem['hFE5D]=8'h84; mem['hFE5E]=8'h27; mem['hFE5F]=8'h0E;
    mem['hFE60]=8'h81; mem['hFE61]=8'h81; mem['hFE62]=8'h26; mem['hFE63]=8'hE7;
    mem['hFE64]=8'h9D; mem['hFE65]=8'h7C; mem['hFE66]=8'h81; mem['hFE67]=8'hA0;
    mem['hFE68]=8'h27; mem['hFE69]=8'h04; mem['hFE6A]=8'h81; mem['hFE6B]=8'hA1;
    mem['hFE6C]=8'h26; mem['hFE6D]=8'hDB; mem['hFE6E]=8'h9D; mem['hFE6F]=8'h7C;
    mem['hFE70]=8'h25; mem['hFE71]=8'h04; mem['hFE72]=8'h9D; mem['hFE73]=8'h82;
    mem['hFE74]=8'h20; mem['hFE75]=8'hD7; mem['hFE76]=8'h9E; mem['hFE77]=8'h83;
    mem['hFE78]=8'h34; mem['hFE79]=8'h10; mem['hFE7A]=8'hBD; mem['hFE7B]=8'hE7;
    mem['hFE7C]=8'h14; mem['hFE7D]=8'h9E; mem['hFE7E]=8'h83; mem['hFE7F]=8'hA6;
    mem['hFE80]=8'h82; mem['hFE81]=8'hBD; mem['hFE82]=8'hFF; mem['hFE83]=8'h73;
    mem['hFE84]=8'h25; mem['hFE85]=8'hF9; mem['hFE86]=8'h30; mem['hFE87]=8'h01;
    mem['hFE88]=8'h1F; mem['hFE89]=8'h10; mem['hFE8A]=8'hE0; mem['hFE8B]=8'h61;
    mem['hFE8C]=8'hC0; mem['hFE8D]=8'h05; mem['hFE8E]=8'h27; mem['hFE8F]=8'h20;
    mem['hFE90]=8'h25; mem['hFE91]=8'h0A; mem['hFE92]=8'h33; mem['hFE93]=8'h84;
    mem['hFE94]=8'h50; mem['hFE95]=8'h30; mem['hFE96]=8'h85; mem['hFE97]=8'hBD;
    mem['hFE98]=8'hFD; mem['hFE99]=8'h25; mem['hFE9A]=8'h20; mem['hFE9B]=8'h14;
    mem['hFE9C]=8'h9F; mem['hFE9D]=8'h47; mem['hFE9E]=8'h9E; mem['hFE9F]=8'h1B;
    mem['hFEA0]=8'h9F; mem['hFEA1]=8'h43; mem['hFEA2]=8'h50; mem['hFEA3]=8'h30;
    mem['hFEA4]=8'h85; mem['hFEA5]=8'h9F; mem['hFEA6]=8'h41; mem['hFEA7]=8'h9F;
    mem['hFEA8]=8'h1B; mem['hFEA9]=8'hBD; mem['hFEAA]=8'hE3; mem['hFEAB]=8'hDB;
    mem['hFEAC]=8'h9E; mem['hFEAD]=8'h45; mem['hFEAE]=8'h9F; mem['hFEAF]=8'h83;
    mem['hFEB0]=8'h35; mem['hFEB1]=8'h10; mem['hFEB2]=8'h86; mem['hFEB3]=8'h01;
    mem['hFEB4]=8'hA7; mem['hFEB5]=8'h84; mem['hFEB6]=8'hA7; mem['hFEB7]=8'h02;
    mem['hFEB8]=8'hA7; mem['hFEB9]=8'h04; mem['hFEBA]=8'hD6; mem['hFEBB]=8'h2B;
    mem['hFEBC]=8'h26; mem['hFEBD]=8'h04; mem['hFEBE]=8'hC6; mem['hFEBF]=8'h01;
    mem['hFEC0]=8'h6C; mem['hFEC1]=8'h02; mem['hFEC2]=8'hE7; mem['hFEC3]=8'h01;
    mem['hFEC4]=8'hD6; mem['hFEC5]=8'h2C; mem['hFEC6]=8'h26; mem['hFEC7]=8'h04;
    mem['hFEC8]=8'hC6; mem['hFEC9]=8'h01; mem['hFECA]=8'h6C; mem['hFECB]=8'h04;
    mem['hFECC]=8'hE7; mem['hFECD]=8'h03; mem['hFECE]=8'h9D; mem['hFECF]=8'h82;
    mem['hFED0]=8'h81; mem['hFED1]=8'h2C; mem['hFED2]=8'h27; mem['hFED3]=8'h9A;
    mem['hFED4]=8'h20; mem['hFED5]=8'h9C; mem['hFED6]=8'h9E; mem['hFED7]=8'h19;
    mem['hFED8]=8'h30; mem['hFED9]=8'h1F; mem['hFEDA]=8'h30; mem['hFEDB]=8'h01;
    mem['hFEDC]=8'hEC; mem['hFEDD]=8'h02; mem['hFEDE]=8'hDD; mem['hFEDF]=8'h68;
    mem['hFEE0]=8'hBD; mem['hFEE1]=8'hFD; mem['hFEE2]=8'hE4; mem['hFEE3]=8'h30;
    mem['hFEE4]=8'h03; mem['hFEE5]=8'h30; mem['hFEE6]=8'h01; mem['hFEE7]=8'hA6;
    mem['hFEE8]=8'h84; mem['hFEE9]=8'h27; mem['hFEEA]=8'hEF; mem['hFEEB]=8'h4A;
    mem['hFEEC]=8'h27; mem['hFEED]=8'h1B; mem['hFEEE]=8'h80; mem['hFEEF]=8'h02;
    mem['hFEF0]=8'h26; mem['hFEF1]=8'hF3; mem['hFEF2]=8'h34; mem['hFEF3]=8'h10;
    mem['hFEF4]=8'h8E; mem['hFEF5]=8'hFF; mem['hFEF6]=8'h33; mem['hFEF7]=8'hBD;
    mem['hFEF8]=8'hF0; mem['hFEF9]=8'hE2; mem['hFEFA]=8'hAE; mem['hFEFB]=8'hE4;
    mem['hFEFC]=8'hEC; mem['hFEFD]=8'h01; mem['hFEFE]=8'hBD; mem['hFEFF]=8'hF5;
    mem['hFF00]=8'h12; mem['hFF01]=8'hBD; mem['hFF02]=8'hF5; mem['hFF03]=8'h0B;
    mem['hFF04]=8'hBD; mem['hFF05]=8'hF0; mem['hFF06]=8'hA2; mem['hFF07]=8'h35;
    mem['hFF08]=8'h10; mem['hFF09]=8'h34; mem['hFF0A]=8'h10; mem['hFF0B]=8'hEC;
    mem['hFF0C]=8'h01; mem['hFF0D]=8'hDD; mem['hFF0E]=8'h52; mem['hFF0F]=8'hBD;
    mem['hFF10]=8'hFB; mem['hFF11]=8'hBE; mem['hFF12]=8'hBD; mem['hFF13]=8'hF5;
    mem['hFF14]=8'h1F; mem['hFF15]=8'h35; mem['hFF16]=8'h40; mem['hFF17]=8'hC6;
    mem['hFF18]=8'h05; mem['hFF19]=8'h30; mem['hFF1A]=8'h01; mem['hFF1B]=8'hA6;
    mem['hFF1C]=8'h84; mem['hFF1D]=8'h27; mem['hFF1E]=8'h05; mem['hFF1F]=8'h5A;
    mem['hFF20]=8'hA7; mem['hFF21]=8'hC0; mem['hFF22]=8'h20; mem['hFF23]=8'hF5;
    mem['hFF24]=8'h30; mem['hFF25]=8'hC4; mem['hFF26]=8'h5D; mem['hFF27]=8'h27;
    mem['hFF28]=8'hBE; mem['hFF29]=8'h31; mem['hFF2A]=8'hC4; mem['hFF2B]=8'h33;
    mem['hFF2C]=8'hC5; mem['hFF2D]=8'hBD; mem['hFF2E]=8'hFD; mem['hFF2F]=8'h25;
    mem['hFF30]=8'h30; mem['hFF31]=8'hA4; mem['hFF32]=8'h20; mem['hFF33]=8'hB3;
    mem['hFF34]=8'h55; mem['hFF35]=8'h4C; mem['hFF36]=8'h20; mem['hFF37]=8'h00;
    mem['hFF38]=8'hBD; mem['hFF39]=8'hEE; mem['hFF3A]=8'hC4; mem['hFF3B]=8'h8E;
    mem['hFF3C]=8'h01; mem['hFF3D]=8'hF0; mem['hFF3E]=8'hC6; mem['hFF3F]=8'h04;
    mem['hFF40]=8'h34; mem['hFF41]=8'h04; mem['hFF42]=8'h5F; mem['hFF43]=8'h86;
    mem['hFF44]=8'h04; mem['hFF45]=8'h08; mem['hFF46]=8'h53; mem['hFF47]=8'h09;
    mem['hFF48]=8'h52; mem['hFF49]=8'h59; mem['hFF4A]=8'h4A; mem['hFF4B]=8'h26;
    mem['hFF4C]=8'hF8; mem['hFF4D]=8'h5D; mem['hFF4E]=8'h26; mem['hFF4F]=8'h0A;
    mem['hFF50]=8'hA6; mem['hFF51]=8'hE4; mem['hFF52]=8'h4A; mem['hFF53]=8'h27;
    mem['hFF54]=8'h05; mem['hFF55]=8'h8C; mem['hFF56]=8'h01; mem['hFF57]=8'hF0;
    mem['hFF58]=8'h27; mem['hFF59]=8'h0C; mem['hFF5A]=8'hCB; mem['hFF5B]=8'h30;
    mem['hFF5C]=8'hC1; mem['hFF5D]=8'h39; mem['hFF5E]=8'h23; mem['hFF5F]=8'h02;
    mem['hFF60]=8'hCB; mem['hFF61]=8'h07; mem['hFF62]=8'hE7; mem['hFF63]=8'h80;
    mem['hFF64]=8'h6F; mem['hFF65]=8'h84; mem['hFF66]=8'h35; mem['hFF67]=8'h04;
    mem['hFF68]=8'h5A; mem['hFF69]=8'h26; mem['hFF6A]=8'hD5; mem['hFF6B]=8'h32;
    mem['hFF6C]=8'h62; mem['hFF6D]=8'h8E; mem['hFF6E]=8'h01; mem['hFF6F]=8'hEF;
    mem['hFF70]=8'h7E; mem['hFF71]=8'hEC; mem['hFF72]=8'h9C; mem['hFF73]=8'h81;
    mem['hFF74]=8'h30; mem['hFF75]=8'h25; mem['hFF76]=8'h04; mem['hFF77]=8'h80;
    mem['hFF78]=8'h3A; mem['hFF79]=8'h80; mem['hFF7A]=8'hC6; mem['hFF7B]=8'h39;
    mem['hFF7C]=8'h81; mem['hFF7D]=8'h89; mem['hFF7E]=8'h10; mem['hFF7F]=8'h27;
    mem['hFF80]=8'hFD; mem['hFF81]=8'hAB; mem['hFF82]=8'h7E; mem['hFF83]=8'hEA;
    mem['hFF84]=8'h00; mem['hFF85]=8'h00; mem['hFF86]=8'h00; mem['hFF87]=8'h00;
    mem['hFF88]=8'h00; mem['hFF89]=8'h00; mem['hFF8A]=8'h00; mem['hFF8B]=8'h00;
    mem['hFF8C]=8'h00; mem['hFF8D]=8'h00; mem['hFF8E]=8'h00; mem['hFF8F]=8'h00;
    mem['hFF90]=8'h00; mem['hFF91]=8'h00; mem['hFF92]=8'h00; mem['hFF93]=8'h00;
    mem['hFF94]=8'h00; mem['hFF95]=8'h00; mem['hFF96]=8'h00; mem['hFF97]=8'h00;
    mem['hFF98]=8'h00; mem['hFF99]=8'h00; mem['hFF9A]=8'h00; mem['hFF9B]=8'h00;
    mem['hFF9C]=8'h00; mem['hFF9D]=8'h00; mem['hFF9E]=8'h00; mem['hFF9F]=8'h00;
    mem['hFFA0]=8'h00; mem['hFFA1]=8'h00; mem['hFFA2]=8'h00; mem['hFFA3]=8'h00;
    mem['hFFA4]=8'h00; mem['hFFA5]=8'h00; mem['hFFA6]=8'h00; mem['hFFA7]=8'h00;
    mem['hFFA8]=8'h00; mem['hFFA9]=8'h00; mem['hFFAA]=8'h00; mem['hFFAB]=8'h00;
    mem['hFFAC]=8'h00; mem['hFFAD]=8'h00; mem['hFFAE]=8'h00; mem['hFFAF]=8'h00;
    mem['hFFB0]=8'h00; mem['hFFB1]=8'h00; mem['hFFB2]=8'h00; mem['hFFB3]=8'h00;
    mem['hFFB4]=8'h00; mem['hFFB5]=8'h00; mem['hFFB6]=8'h00; mem['hFFB7]=8'h00;
    mem['hFFB8]=8'h00; mem['hFFB9]=8'h00; mem['hFFBA]=8'h00; mem['hFFBB]=8'h00;
    mem['hFFBC]=8'h00; mem['hFFBD]=8'h00; mem['hFFBE]=8'h00; mem['hFFBF]=8'h00;
    mem['hFFC0]=8'h00; mem['hFFC1]=8'h00; mem['hFFC2]=8'h00; mem['hFFC3]=8'h00;
    mem['hFFC4]=8'h00; mem['hFFC5]=8'h00; mem['hFFC6]=8'h00; mem['hFFC7]=8'h00;
    mem['hFFC8]=8'h00; mem['hFFC9]=8'h00; mem['hFFCA]=8'h00; mem['hFFCB]=8'h00;
    mem['hFFCC]=8'h00; mem['hFFCD]=8'h00; mem['hFFCE]=8'h00; mem['hFFCF]=8'h00;
    mem['hFFD0]=8'h00; mem['hFFD1]=8'h00; mem['hFFD2]=8'h00; mem['hFFD3]=8'h00;
    mem['hFFD4]=8'h00; mem['hFFD5]=8'h00; mem['hFFD6]=8'h00; mem['hFFD7]=8'h00;
    mem['hFFD8]=8'h00; mem['hFFD9]=8'h00; mem['hFFDA]=8'h00; mem['hFFDB]=8'h00;
    mem['hFFDC]=8'h00; mem['hFFDD]=8'h00; mem['hFFDE]=8'h00; mem['hFFDF]=8'h00;
    mem['hFFE0]=8'h00; mem['hFFE1]=8'h00; mem['hFFE2]=8'h00; mem['hFFE3]=8'h00;
    mem['hFFE4]=8'h00; mem['hFFE5]=8'h00; mem['hFFE6]=8'h00; mem['hFFE7]=8'h00;
    mem['hFFE8]=8'h00; mem['hFFE9]=8'h00; mem['hFFEA]=8'h00; mem['hFFEB]=8'h00;
    mem['hFFEC]=8'h00; mem['hFFED]=8'h00; mem['hFFEE]=8'h00; mem['hFFEF]=8'h00;
    mem['hFFF0]=8'h00; mem['hFFF1]=8'h00; mem['hFFF2]=8'h00; mem['hFFF3]=8'h9B;
    mem['hFFF4]=8'h00; mem['hFFF5]=8'h9E; mem['hFFF6]=8'h00; mem['hFFF7]=8'hAA;
    mem['hFFF8]=8'h00; mem['hFFF9]=8'hA7; mem['hFFFA]=8'h00; mem['hFFFB]=8'hA1;
    mem['hFFFC]=8'h00; mem['hFFFD]=8'hA4; mem['hFFFE]=8'hE0; mem['hFFFF]=8'h46;
end
