// rom.v
// to be included from the top module at the comple

initial
begin
    mem['h0000]=8'hF3; mem['h0001]=8'h31; mem['h0002]=8'hED; mem['h0003]=8'h80;
    mem['h0004]=8'hC3; mem['h0005]=8'h1B; mem['h0006]=8'h00; mem['h0007]=8'hFF;
    mem['h0008]=8'hC3; mem['h0009]=8'hC9; mem['h000A]=8'h00; mem['h000B]=8'hFF;
    mem['h000C]=8'hFF; mem['h000D]=8'hFF; mem['h000E]=8'hFF; mem['h000F]=8'hFF;
    mem['h0010]=8'hC3; mem['h0011]=8'h9D; mem['h0012]=8'h00; mem['h0013]=8'hFF;
    mem['h0014]=8'hFF; mem['h0015]=8'hFF; mem['h0016]=8'hFF; mem['h0017]=8'hFF;
    mem['h0018]=8'hC3; mem['h0019]=8'hC3; mem['h001A]=8'h00; mem['h001B]=8'h21;
    mem['h001C]=8'h00; mem['h001D]=8'h80; mem['h001E]=8'h11; mem['h001F]=8'h00;
    mem['h0020]=8'h80; mem['h0021]=8'h01; mem['h0022]=8'h00; mem['h0023]=8'h40;
    mem['h0024]=8'hED; mem['h0025]=8'hB0; mem['h0026]=8'hAF; mem['h0027]=8'h32;
    mem['h0028]=8'h00; mem['h0029]=8'h80; mem['h002A]=8'h32; mem['h002B]=8'h01;
    mem['h002C]=8'h80; mem['h002D]=8'h32; mem['h002E]=8'h02; mem['h002F]=8'h80;
    mem['h0030]=8'hED; mem['h0031]=8'h5E; mem['h0032]=8'h21; mem['h0033]=8'h60;
    mem['h0034]=8'h00; mem['h0035]=8'h7C; mem['h0036]=8'hED; mem['h0037]=8'h47;
    mem['h0038]=8'h21; mem['h0039]=8'h4E; mem['h003A]=8'h00; mem['h003B]=8'h0E;
    mem['h003C]=8'h01; mem['h003D]=8'h06; mem['h003E]=8'h09; mem['h003F]=8'hED;
    mem['h0040]=8'hB3; mem['h0041]=8'h21; mem['h0042]=8'h57; mem['h0043]=8'h00;
    mem['h0044]=8'h0E; mem['h0045]=8'h03; mem['h0046]=8'h06; mem['h0047]=8'h05;
    mem['h0048]=8'hED; mem['h0049]=8'hB3; mem['h004A]=8'hFB; mem['h004B]=8'hC3;
    mem['h004C]=8'hD4; mem['h004D]=8'h00; mem['h004E]=8'h18; mem['h004F]=8'h01;
    mem['h0050]=8'h14; mem['h0051]=8'h04; mem['h0052]=8'h44; mem['h0053]=8'h05;
    mem['h0054]=8'hEA; mem['h0055]=8'h03; mem['h0056]=8'hC1; mem['h0057]=8'h18;
    mem['h0058]=8'h01; mem['h0059]=8'h04; mem['h005A]=8'h02; mem['h005B]=8'h60;
    mem['h005C]=8'hFF; mem['h005D]=8'hFF; mem['h005E]=8'hFF; mem['h005F]=8'hFF;
    mem['h0060]=8'h00; mem['h0061]=8'h00; mem['h0062]=8'h00; mem['h0063]=8'h00;
    mem['h0064]=8'h00; mem['h0065]=8'h00; mem['h0066]=8'h00; mem['h0067]=8'h00;
    mem['h0068]=8'h70; mem['h0069]=8'h00; mem['h006A]=8'h70; mem['h006B]=8'h00;
    mem['h006C]=8'h73; mem['h006D]=8'h00; mem['h006E]=8'h70; mem['h006F]=8'h00;
    mem['h0070]=8'hFB; mem['h0071]=8'hED; mem['h0072]=8'h4D; mem['h0073]=8'hF5;
    mem['h0074]=8'hC5; mem['h0075]=8'hD5; mem['h0076]=8'hE5; mem['h0077]=8'hDB;
    mem['h0078]=8'h00; mem['h0079]=8'h57; mem['h007A]=8'h3A; mem['h007B]=8'h00;
    mem['h007C]=8'h80; mem['h007D]=8'hFE; mem['h007E]=8'h40; mem['h007F]=8'h28;
    mem['h0080]=8'h15; mem['h0081]=8'h3C; mem['h0082]=8'h32; mem['h0083]=8'h00;
    mem['h0084]=8'h80; mem['h0085]=8'h3A; mem['h0086]=8'h02; mem['h0087]=8'h80;
    mem['h0088]=8'h4F; mem['h0089]=8'h06; mem['h008A]=8'h00; mem['h008B]=8'h21;
    mem['h008C]=8'h03; mem['h008D]=8'h80; mem['h008E]=8'h09; mem['h008F]=8'h72;
    mem['h0090]=8'h3C; mem['h0091]=8'hE6; mem['h0092]=8'h3F; mem['h0093]=8'h32;
    mem['h0094]=8'h02; mem['h0095]=8'h80; mem['h0096]=8'hE1; mem['h0097]=8'hD1;
    mem['h0098]=8'hC1; mem['h0099]=8'hF1; mem['h009A]=8'hFB; mem['h009B]=8'hED;
    mem['h009C]=8'h4D; mem['h009D]=8'hC5; mem['h009E]=8'hD5; mem['h009F]=8'hE5;
    mem['h00A0]=8'h3A; mem['h00A1]=8'h00; mem['h00A2]=8'h80; mem['h00A3]=8'hFE;
    mem['h00A4]=8'h00; mem['h00A5]=8'h28; mem['h00A6]=8'hF9; mem['h00A7]=8'hF3;
    mem['h00A8]=8'h3D; mem['h00A9]=8'h32; mem['h00AA]=8'h00; mem['h00AB]=8'h80;
    mem['h00AC]=8'h3A; mem['h00AD]=8'h01; mem['h00AE]=8'h80; mem['h00AF]=8'h4F;
    mem['h00B0]=8'h06; mem['h00B1]=8'h00; mem['h00B2]=8'h21; mem['h00B3]=8'h03;
    mem['h00B4]=8'h80; mem['h00B5]=8'h09; mem['h00B6]=8'h56; mem['h00B7]=8'h3C;
    mem['h00B8]=8'hE6; mem['h00B9]=8'h3F; mem['h00BA]=8'h32; mem['h00BB]=8'h01;
    mem['h00BC]=8'h80; mem['h00BD]=8'h7A; mem['h00BE]=8'hFB; mem['h00BF]=8'hE1;
    mem['h00C0]=8'hD1; mem['h00C1]=8'hC1; mem['h00C2]=8'hC9; mem['h00C3]=8'h3A;
    mem['h00C4]=8'h00; mem['h00C5]=8'h80; mem['h00C6]=8'hFE; mem['h00C7]=8'h00;
    mem['h00C8]=8'hC9; mem['h00C9]=8'hF5; mem['h00CA]=8'hDB; mem['h00CB]=8'h01;
    mem['h00CC]=8'hCB; mem['h00CD]=8'h57; mem['h00CE]=8'h28; mem['h00CF]=8'hFA;
    mem['h00D0]=8'hF1; mem['h00D1]=8'hD3; mem['h00D2]=8'h00; mem['h00D3]=8'hC9;
    mem['h00D4]=8'hC3; mem['h00D5]=8'hDA; mem['h00D6]=8'h00; mem['h00D7]=8'hC3;
    mem['h00D8]=8'h4F; mem['h00D9]=8'h01; mem['h00DA]=8'hC3; mem['h00DB]=8'hE1;
    mem['h00DC]=8'h00; mem['h00DD]=8'h92; mem['h00DE]=8'h09; mem['h00DF]=8'h08;
    mem['h00E0]=8'h11; mem['h00E1]=8'h21; mem['h00E2]=8'h45; mem['h00E3]=8'h80;
    mem['h00E4]=8'hF9; mem['h00E5]=8'hC3; mem['h00E6]=8'h23; mem['h00E7]=8'h1D;
    mem['h00E8]=8'h11; mem['h00E9]=8'hB9; mem['h00EA]=8'h03; mem['h00EB]=8'h06;
    mem['h00EC]=8'h63; mem['h00ED]=8'h21; mem['h00EE]=8'h45; mem['h00EF]=8'h80;
    mem['h00F0]=8'h1A; mem['h00F1]=8'h77; mem['h00F2]=8'h23; mem['h00F3]=8'h13;
    mem['h00F4]=8'h05; mem['h00F5]=8'hC2; mem['h00F6]=8'hF0; mem['h00F7]=8'h00;
    mem['h00F8]=8'hF9; mem['h00F9]=8'hCD; mem['h00FA]=8'hBA; mem['h00FB]=8'h05;
    mem['h00FC]=8'hCD; mem['h00FD]=8'h88; mem['h00FE]=8'h0B; mem['h00FF]=8'h32;
    mem['h0100]=8'hEF; mem['h0101]=8'h80; mem['h0102]=8'h32; mem['h0103]=8'h3E;
    mem['h0104]=8'h81; mem['h0105]=8'h21; mem['h0106]=8'hA2; mem['h0107]=8'h81;
    mem['h0108]=8'h23; mem['h0109]=8'h7C; mem['h010A]=8'hB5; mem['h010B]=8'hCA;
    mem['h010C]=8'h17; mem['h010D]=8'h01; mem['h010E]=8'h7E; mem['h010F]=8'h47;
    mem['h0110]=8'h2F; mem['h0111]=8'h77; mem['h0112]=8'hBE; mem['h0113]=8'h70;
    mem['h0114]=8'hCA; mem['h0115]=8'h08; mem['h0116]=8'h01; mem['h0117]=8'h2B;
    mem['h0118]=8'h11; mem['h0119]=8'hA1; mem['h011A]=8'h81; mem['h011B]=8'hCD;
    mem['h011C]=8'h50; mem['h011D]=8'h07; mem['h011E]=8'hDA; mem['h011F]=8'h58;
    mem['h0120]=8'h01; mem['h0121]=8'h11; mem['h0122]=8'hCE; mem['h0123]=8'hFF;
    mem['h0124]=8'h22; mem['h0125]=8'hF4; mem['h0126]=8'h80; mem['h0127]=8'h19;
    mem['h0128]=8'h22; mem['h0129]=8'h9F; mem['h012A]=8'h80; mem['h012B]=8'hCD;
    mem['h012C]=8'h95; mem['h012D]=8'h05; mem['h012E]=8'h2A; mem['h012F]=8'h9F;
    mem['h0130]=8'h80; mem['h0131]=8'h11; mem['h0132]=8'hEF; mem['h0133]=8'hFF;
    mem['h0134]=8'h19; mem['h0135]=8'h11; mem['h0136]=8'h3E; mem['h0137]=8'h81;
    mem['h0138]=8'h7D; mem['h0139]=8'h93; mem['h013A]=8'h6F; mem['h013B]=8'h7C;
    mem['h013C]=8'h9A; mem['h013D]=8'h67; mem['h013E]=8'hE5; mem['h013F]=8'h21;
    mem['h0140]=8'h70; mem['h0141]=8'h01; mem['h0142]=8'hCD; mem['h0143]=8'h26;
    mem['h0144]=8'h12; mem['h0145]=8'hE1; mem['h0146]=8'hCD; mem['h0147]=8'hC9;
    mem['h0148]=8'h18; mem['h0149]=8'h21; mem['h014A]=8'h61; mem['h014B]=8'h01;
    mem['h014C]=8'hCD; mem['h014D]=8'h26; mem['h014E]=8'h12; mem['h014F]=8'h31;
    mem['h0150]=8'hAB; mem['h0151]=8'h80; mem['h0152]=8'hCD; mem['h0153]=8'hBA;
    mem['h0154]=8'h05; mem['h0155]=8'hC3; mem['h0156]=8'hD3; mem['h0157]=8'h04;
    mem['h0158]=8'h21; mem['h0159]=8'hA7; mem['h015A]=8'h01; mem['h015B]=8'hCD;
    mem['h015C]=8'h26; mem['h015D]=8'h12; mem['h015E]=8'hC3; mem['h015F]=8'h5E;
    mem['h0160]=8'h01; mem['h0161]=8'h20; mem['h0162]=8'h42; mem['h0163]=8'h79;
    mem['h0164]=8'h74; mem['h0165]=8'h65; mem['h0166]=8'h73; mem['h0167]=8'h20;
    mem['h0168]=8'h66; mem['h0169]=8'h72; mem['h016A]=8'h65; mem['h016B]=8'h65;
    mem['h016C]=8'h0D; mem['h016D]=8'h0A; mem['h016E]=8'h00; mem['h016F]=8'h00;
    mem['h0170]=8'h5A; mem['h0171]=8'h38; mem['h0172]=8'h30; mem['h0173]=8'h20;
    mem['h0174]=8'h42; mem['h0175]=8'h41; mem['h0176]=8'h53; mem['h0177]=8'h49;
    mem['h0178]=8'h43; mem['h0179]=8'h20; mem['h017A]=8'h56; mem['h017B]=8'h65;
    mem['h017C]=8'h72; mem['h017D]=8'h20; mem['h017E]=8'h34; mem['h017F]=8'h2E;
    mem['h0180]=8'h37; mem['h0181]=8'h62; mem['h0182]=8'h0D; mem['h0183]=8'h0A;
    mem['h0184]=8'h43; mem['h0185]=8'h6F; mem['h0186]=8'h70; mem['h0187]=8'h79;
    mem['h0188]=8'h72; mem['h0189]=8'h69; mem['h018A]=8'h67; mem['h018B]=8'h68;
    mem['h018C]=8'h74; mem['h018D]=8'h20; mem['h018E]=8'h28; mem['h018F]=8'h43;
    mem['h0190]=8'h29; mem['h0191]=8'h20; mem['h0192]=8'h31; mem['h0193]=8'h39;
    mem['h0194]=8'h37; mem['h0195]=8'h38; mem['h0196]=8'h20; mem['h0197]=8'h62;
    mem['h0198]=8'h79; mem['h0199]=8'h20; mem['h019A]=8'h4D; mem['h019B]=8'h69;
    mem['h019C]=8'h63; mem['h019D]=8'h72; mem['h019E]=8'h6F; mem['h019F]=8'h73;
    mem['h01A0]=8'h6F; mem['h01A1]=8'h66; mem['h01A2]=8'h74; mem['h01A3]=8'h0D;
    mem['h01A4]=8'h0A; mem['h01A5]=8'h00; mem['h01A6]=8'h00; mem['h01A7]=8'h4D;
    mem['h01A8]=8'h65; mem['h01A9]=8'h6D; mem['h01AA]=8'h6F; mem['h01AB]=8'h72;
    mem['h01AC]=8'h79; mem['h01AD]=8'h20; mem['h01AE]=8'h73; mem['h01AF]=8'h69;
    mem['h01B0]=8'h7A; mem['h01B1]=8'h65; mem['h01B2]=8'h20; mem['h01B3]=8'h6E;
    mem['h01B4]=8'h6F; mem['h01B5]=8'h74; mem['h01B6]=8'h20; mem['h01B7]=8'h65;
    mem['h01B8]=8'h6E; mem['h01B9]=8'h6F; mem['h01BA]=8'h75; mem['h01BB]=8'h67;
    mem['h01BC]=8'h68; mem['h01BD]=8'h0D; mem['h01BE]=8'h0A; mem['h01BF]=8'h54;
    mem['h01C0]=8'h68; mem['h01C1]=8'h65; mem['h01C2]=8'h20; mem['h01C3]=8'h73;
    mem['h01C4]=8'h79; mem['h01C5]=8'h73; mem['h01C6]=8'h74; mem['h01C7]=8'h65;
    mem['h01C8]=8'h6D; mem['h01C9]=8'h20; mem['h01CA]=8'h69; mem['h01CB]=8'h73;
    mem['h01CC]=8'h20; mem['h01CD]=8'h73; mem['h01CE]=8'h74; mem['h01CF]=8'h6F;
    mem['h01D0]=8'h70; mem['h01D1]=8'h70; mem['h01D2]=8'h65; mem['h01D3]=8'h64;
    mem['h01D4]=8'h2E; mem['h01D5]=8'h0D; mem['h01D6]=8'h0A; mem['h01D7]=8'h00;
    mem['h01D8]=8'h00; mem['h01D9]=8'h3E; mem['h01DA]=8'h17; mem['h01DB]=8'h02;
    mem['h01DC]=8'h18; mem['h01DD]=8'h54; mem['h01DE]=8'h17; mem['h01DF]=8'h48;
    mem['h01E0]=8'h80; mem['h01E1]=8'hE6; mem['h01E2]=8'h10; mem['h01E3]=8'h6B;
    mem['h01E4]=8'h14; mem['h01E5]=8'h14; mem['h01E6]=8'h11; mem['h01E7]=8'hC8;
    mem['h01E8]=8'h19; mem['h01E9]=8'hA7; mem['h01EA]=8'h1A; mem['h01EB]=8'hE3;
    mem['h01EC]=8'h15; mem['h01ED]=8'h16; mem['h01EE]=8'h1A; mem['h01EF]=8'h1C;
    mem['h01F0]=8'h1B; mem['h01F1]=8'h22; mem['h01F2]=8'h1B; mem['h01F3]=8'h83;
    mem['h01F4]=8'h1B; mem['h01F5]=8'h98; mem['h01F6]=8'h1B; mem['h01F7]=8'hBF;
    mem['h01F8]=8'h14; mem['h01F9]=8'h03; mem['h01FA]=8'h1C; mem['h01FB]=8'h96;
    mem['h01FC]=8'h80; mem['h01FD]=8'h98; mem['h01FE]=8'h13; mem['h01FF]=8'hB0;
    mem['h0200]=8'h11; mem['h0201]=8'h32; mem['h0202]=8'h14; mem['h0203]=8'hA7;
    mem['h0204]=8'h13; mem['h0205]=8'hB8; mem['h0206]=8'h13; mem['h0207]=8'h25;
    mem['h0208]=8'h1C; mem['h0209]=8'hB8; mem['h020A]=8'h1C; mem['h020B]=8'hC8;
    mem['h020C]=8'h13; mem['h020D]=8'hF8; mem['h020E]=8'h13; mem['h020F]=8'h02;
    mem['h0210]=8'h14; mem['h0211]=8'hC5; mem['h0212]=8'h4E; mem['h0213]=8'h44;
    mem['h0214]=8'hC6; mem['h0215]=8'h4F; mem['h0216]=8'h52; mem['h0217]=8'hCE;
    mem['h0218]=8'h45; mem['h0219]=8'h58; mem['h021A]=8'h54; mem['h021B]=8'hC4;
    mem['h021C]=8'h41; mem['h021D]=8'h54; mem['h021E]=8'h41; mem['h021F]=8'hC9;
    mem['h0220]=8'h4E; mem['h0221]=8'h50; mem['h0222]=8'h55; mem['h0223]=8'h54;
    mem['h0224]=8'hC4; mem['h0225]=8'h49; mem['h0226]=8'h4D; mem['h0227]=8'hD2;
    mem['h0228]=8'h45; mem['h0229]=8'h41; mem['h022A]=8'h44; mem['h022B]=8'hCC;
    mem['h022C]=8'h45; mem['h022D]=8'h54; mem['h022E]=8'hC7; mem['h022F]=8'h4F;
    mem['h0230]=8'h54; mem['h0231]=8'h4F; mem['h0232]=8'hD2; mem['h0233]=8'h55;
    mem['h0234]=8'h4E; mem['h0235]=8'hC9; mem['h0236]=8'h46; mem['h0237]=8'hD2;
    mem['h0238]=8'h45; mem['h0239]=8'h53; mem['h023A]=8'h54; mem['h023B]=8'h4F;
    mem['h023C]=8'h52; mem['h023D]=8'h45; mem['h023E]=8'hC7; mem['h023F]=8'h4F;
    mem['h0240]=8'h53; mem['h0241]=8'h55; mem['h0242]=8'h42; mem['h0243]=8'hD2;
    mem['h0244]=8'h45; mem['h0245]=8'h54; mem['h0246]=8'h55; mem['h0247]=8'h52;
    mem['h0248]=8'h4E; mem['h0249]=8'hD2; mem['h024A]=8'h45; mem['h024B]=8'h4D;
    mem['h024C]=8'hD3; mem['h024D]=8'h54; mem['h024E]=8'h4F; mem['h024F]=8'h50;
    mem['h0250]=8'hCF; mem['h0251]=8'h55; mem['h0252]=8'h54; mem['h0253]=8'hCF;
    mem['h0254]=8'h4E; mem['h0255]=8'hCE; mem['h0256]=8'h55; mem['h0257]=8'h4C;
    mem['h0258]=8'h4C; mem['h0259]=8'hD7; mem['h025A]=8'h41; mem['h025B]=8'h49;
    mem['h025C]=8'h54; mem['h025D]=8'hC4; mem['h025E]=8'h45; mem['h025F]=8'h46;
    mem['h0260]=8'hD0; mem['h0261]=8'h4F; mem['h0262]=8'h4B; mem['h0263]=8'h45;
    mem['h0264]=8'hC4; mem['h0265]=8'h4F; mem['h0266]=8'h4B; mem['h0267]=8'h45;
    mem['h0268]=8'hD3; mem['h0269]=8'h43; mem['h026A]=8'h52; mem['h026B]=8'h45;
    mem['h026C]=8'h45; mem['h026D]=8'h4E; mem['h026E]=8'hCC; mem['h026F]=8'h49;
    mem['h0270]=8'h4E; mem['h0271]=8'h45; mem['h0272]=8'h53; mem['h0273]=8'hC3;
    mem['h0274]=8'h4C; mem['h0275]=8'h53; mem['h0276]=8'hD7; mem['h0277]=8'h49;
    mem['h0278]=8'h44; mem['h0279]=8'h54; mem['h027A]=8'h48; mem['h027B]=8'hCD;
    mem['h027C]=8'h4F; mem['h027D]=8'h4E; mem['h027E]=8'h49; mem['h027F]=8'h54;
    mem['h0280]=8'h4F; mem['h0281]=8'h52; mem['h0282]=8'hD3; mem['h0283]=8'h45;
    mem['h0284]=8'h54; mem['h0285]=8'hD2; mem['h0286]=8'h45; mem['h0287]=8'h53;
    mem['h0288]=8'h45; mem['h0289]=8'h54; mem['h028A]=8'hD0; mem['h028B]=8'h52;
    mem['h028C]=8'h49; mem['h028D]=8'h4E; mem['h028E]=8'h54; mem['h028F]=8'hC3;
    mem['h0290]=8'h4F; mem['h0291]=8'h4E; mem['h0292]=8'h54; mem['h0293]=8'hCC;
    mem['h0294]=8'h49; mem['h0295]=8'h53; mem['h0296]=8'h54; mem['h0297]=8'hC3;
    mem['h0298]=8'h4C; mem['h0299]=8'h45; mem['h029A]=8'h41; mem['h029B]=8'h52;
    mem['h029C]=8'hC3; mem['h029D]=8'h4C; mem['h029E]=8'h4F; mem['h029F]=8'h41;
    mem['h02A0]=8'h44; mem['h02A1]=8'hC3; mem['h02A2]=8'h53; mem['h02A3]=8'h41;
    mem['h02A4]=8'h56; mem['h02A5]=8'h45; mem['h02A6]=8'hCE; mem['h02A7]=8'h45;
    mem['h02A8]=8'h57; mem['h02A9]=8'hD4; mem['h02AA]=8'h41; mem['h02AB]=8'h42;
    mem['h02AC]=8'h28; mem['h02AD]=8'hD4; mem['h02AE]=8'h4F; mem['h02AF]=8'hC6;
    mem['h02B0]=8'h4E; mem['h02B1]=8'hD3; mem['h02B2]=8'h50; mem['h02B3]=8'h43;
    mem['h02B4]=8'h28; mem['h02B5]=8'hD4; mem['h02B6]=8'h48; mem['h02B7]=8'h45;
    mem['h02B8]=8'h4E; mem['h02B9]=8'hCE; mem['h02BA]=8'h4F; mem['h02BB]=8'h54;
    mem['h02BC]=8'hD3; mem['h02BD]=8'h54; mem['h02BE]=8'h45; mem['h02BF]=8'h50;
    mem['h02C0]=8'hAB; mem['h02C1]=8'hAD; mem['h02C2]=8'hAA; mem['h02C3]=8'hAF;
    mem['h02C4]=8'hDE; mem['h02C5]=8'hC1; mem['h02C6]=8'h4E; mem['h02C7]=8'h44;
    mem['h02C8]=8'hCF; mem['h02C9]=8'h52; mem['h02CA]=8'hBE; mem['h02CB]=8'hBD;
    mem['h02CC]=8'hBC; mem['h02CD]=8'hD3; mem['h02CE]=8'h47; mem['h02CF]=8'h4E;
    mem['h02D0]=8'hC9; mem['h02D1]=8'h4E; mem['h02D2]=8'h54; mem['h02D3]=8'hC1;
    mem['h02D4]=8'h42; mem['h02D5]=8'h53; mem['h02D6]=8'hD5; mem['h02D7]=8'h53;
    mem['h02D8]=8'h52; mem['h02D9]=8'hC6; mem['h02DA]=8'h52; mem['h02DB]=8'h45;
    mem['h02DC]=8'hC9; mem['h02DD]=8'h4E; mem['h02DE]=8'h50; mem['h02DF]=8'hD0;
    mem['h02E0]=8'h4F; mem['h02E1]=8'h53; mem['h02E2]=8'hD3; mem['h02E3]=8'h51;
    mem['h02E4]=8'h52; mem['h02E5]=8'hD2; mem['h02E6]=8'h4E; mem['h02E7]=8'h44;
    mem['h02E8]=8'hCC; mem['h02E9]=8'h4F; mem['h02EA]=8'h47; mem['h02EB]=8'hC5;
    mem['h02EC]=8'h58; mem['h02ED]=8'h50; mem['h02EE]=8'hC3; mem['h02EF]=8'h4F;
    mem['h02F0]=8'h53; mem['h02F1]=8'hD3; mem['h02F2]=8'h49; mem['h02F3]=8'h4E;
    mem['h02F4]=8'hD4; mem['h02F5]=8'h41; mem['h02F6]=8'h4E; mem['h02F7]=8'hC1;
    mem['h02F8]=8'h54; mem['h02F9]=8'h4E; mem['h02FA]=8'hD0; mem['h02FB]=8'h45;
    mem['h02FC]=8'h45; mem['h02FD]=8'h4B; mem['h02FE]=8'hC4; mem['h02FF]=8'h45;
    mem['h0300]=8'h45; mem['h0301]=8'h4B; mem['h0302]=8'hD0; mem['h0303]=8'h4F;
    mem['h0304]=8'h49; mem['h0305]=8'h4E; mem['h0306]=8'h54; mem['h0307]=8'hCC;
    mem['h0308]=8'h45; mem['h0309]=8'h4E; mem['h030A]=8'hD3; mem['h030B]=8'h54;
    mem['h030C]=8'h52; mem['h030D]=8'h24; mem['h030E]=8'hD6; mem['h030F]=8'h41;
    mem['h0310]=8'h4C; mem['h0311]=8'hC1; mem['h0312]=8'h53; mem['h0313]=8'h43;
    mem['h0314]=8'hC3; mem['h0315]=8'h48; mem['h0316]=8'h52; mem['h0317]=8'h24;
    mem['h0318]=8'hC8; mem['h0319]=8'h45; mem['h031A]=8'h58; mem['h031B]=8'h24;
    mem['h031C]=8'hC2; mem['h031D]=8'h49; mem['h031E]=8'h4E; mem['h031F]=8'h24;
    mem['h0320]=8'hCC; mem['h0321]=8'h45; mem['h0322]=8'h46; mem['h0323]=8'h54;
    mem['h0324]=8'h24; mem['h0325]=8'hD2; mem['h0326]=8'h49; mem['h0327]=8'h47;
    mem['h0328]=8'h48; mem['h0329]=8'h54; mem['h032A]=8'h24; mem['h032B]=8'hCD;
    mem['h032C]=8'h49; mem['h032D]=8'h44; mem['h032E]=8'h24; mem['h032F]=8'h80;
    mem['h0330]=8'h2A; mem['h0331]=8'h09; mem['h0332]=8'h27; mem['h0333]=8'h08;
    mem['h0334]=8'h02; mem['h0335]=8'h0D; mem['h0336]=8'h77; mem['h0337]=8'h0A;
    mem['h0338]=8'h09; mem['h0339]=8'h0C; mem['h033A]=8'h3E; mem['h033B]=8'h0F;
    mem['h033C]=8'h38; mem['h033D]=8'h0C; mem['h033E]=8'h8E; mem['h033F]=8'h0A;
    mem['h0340]=8'h34; mem['h0341]=8'h0A; mem['h0342]=8'h17; mem['h0343]=8'h0A;
    mem['h0344]=8'h06; mem['h0345]=8'h0B; mem['h0346]=8'hF0; mem['h0347]=8'h08;
    mem['h0348]=8'h23; mem['h0349]=8'h0A; mem['h034A]=8'h52; mem['h034B]=8'h0A;
    mem['h034C]=8'h79; mem['h034D]=8'h0A; mem['h034E]=8'h28; mem['h034F]=8'h09;
    mem['h0350]=8'h77; mem['h0351]=8'h14; mem['h0352]=8'hE8; mem['h0353]=8'h0A;
    mem['h0354]=8'h69; mem['h0355]=8'h09; mem['h0356]=8'h7D; mem['h0357]=8'h14;
    mem['h0358]=8'h1C; mem['h0359]=8'h11; mem['h035A]=8'hC6; mem['h035B]=8'h14;
    mem['h035C]=8'h0E; mem['h035D]=8'h1C; mem['h035E]=8'h79; mem['h035F]=8'h0A;
    mem['h0360]=8'hF4; mem['h0361]=8'h1B; mem['h0362]=8'hE7; mem['h0363]=8'h1B;
    mem['h0364]=8'hEC; mem['h0365]=8'h1B; mem['h0366]=8'h20; mem['h0367]=8'h1D;
    mem['h0368]=8'h99; mem['h0369]=8'h80; mem['h036A]=8'h9C; mem['h036B]=8'h80;
    mem['h036C]=8'h2A; mem['h036D]=8'h0B; mem['h036E]=8'h56; mem['h036F]=8'h09;
    mem['h0370]=8'h9C; mem['h0371]=8'h07; mem['h0372]=8'hD1; mem['h0373]=8'h09;
    mem['h0374]=8'h79; mem['h0375]=8'h0A; mem['h0376]=8'h79; mem['h0377]=8'h0A;
    mem['h0378]=8'h94; mem['h0379]=8'h05; mem['h037A]=8'h79; mem['h037B]=8'hB0;
    mem['h037C]=8'h18; mem['h037D]=8'h79; mem['h037E]=8'hE4; mem['h037F]=8'h14;
    mem['h0380]=8'h7C; mem['h0381]=8'h22; mem['h0382]=8'h16; mem['h0383]=8'h7C;
    mem['h0384]=8'h83; mem['h0385]=8'h16; mem['h0386]=8'h7F; mem['h0387]=8'hD1;
    mem['h0388]=8'h19; mem['h0389]=8'h50; mem['h038A]=8'h97; mem['h038B]=8'h0E;
    mem['h038C]=8'h46; mem['h038D]=8'h96; mem['h038E]=8'h0E; mem['h038F]=8'h4E;
    mem['h0390]=8'h46; mem['h0391]=8'h53; mem['h0392]=8'h4E; mem['h0393]=8'h52;
    mem['h0394]=8'h47; mem['h0395]=8'h4F; mem['h0396]=8'h44; mem['h0397]=8'h46;
    mem['h0398]=8'h43; mem['h0399]=8'h4F; mem['h039A]=8'h56; mem['h039B]=8'h4F;
    mem['h039C]=8'h4D; mem['h039D]=8'h55; mem['h039E]=8'h4C; mem['h039F]=8'h42;
    mem['h03A0]=8'h53; mem['h03A1]=8'h44; mem['h03A2]=8'h44; mem['h03A3]=8'h2F;
    mem['h03A4]=8'h30; mem['h03A5]=8'h49; mem['h03A6]=8'h44; mem['h03A7]=8'h54;
    mem['h03A8]=8'h4D; mem['h03A9]=8'h4F; mem['h03AA]=8'h53; mem['h03AB]=8'h4C;
    mem['h03AC]=8'h53; mem['h03AD]=8'h53; mem['h03AE]=8'h54; mem['h03AF]=8'h43;
    mem['h03B0]=8'h4E; mem['h03B1]=8'h55; mem['h03B2]=8'h46; mem['h03B3]=8'h4D;
    mem['h03B4]=8'h4F; mem['h03B5]=8'h48; mem['h03B6]=8'h58; mem['h03B7]=8'h42;
    mem['h03B8]=8'h4E; mem['h03B9]=8'hC3; mem['h03BA]=8'h4F; mem['h03BB]=8'h01;
    mem['h03BC]=8'hC3; mem['h03BD]=8'hA7; mem['h03BE]=8'h09; mem['h03BF]=8'hD3;
    mem['h03C0]=8'h00; mem['h03C1]=8'hC9; mem['h03C2]=8'hD6; mem['h03C3]=8'h00;
    mem['h03C4]=8'h6F; mem['h03C5]=8'h7C; mem['h03C6]=8'hDE; mem['h03C7]=8'h00;
    mem['h03C8]=8'h67; mem['h03C9]=8'h78; mem['h03CA]=8'hDE; mem['h03CB]=8'h00;
    mem['h03CC]=8'h47; mem['h03CD]=8'h3E; mem['h03CE]=8'h00; mem['h03CF]=8'hC9;
    mem['h03D0]=8'h00; mem['h03D1]=8'h00; mem['h03D2]=8'h00; mem['h03D3]=8'h35;
    mem['h03D4]=8'h4A; mem['h03D5]=8'hCA; mem['h03D6]=8'h99; mem['h03D7]=8'h39;
    mem['h03D8]=8'h1C; mem['h03D9]=8'h76; mem['h03DA]=8'h98; mem['h03DB]=8'h22;
    mem['h03DC]=8'h95; mem['h03DD]=8'hB3; mem['h03DE]=8'h98; mem['h03DF]=8'h0A;
    mem['h03E0]=8'hDD; mem['h03E1]=8'h47; mem['h03E2]=8'h98; mem['h03E3]=8'h53;
    mem['h03E4]=8'hD1; mem['h03E5]=8'h99; mem['h03E6]=8'h99; mem['h03E7]=8'h0A;
    mem['h03E8]=8'h1A; mem['h03E9]=8'h9F; mem['h03EA]=8'h98; mem['h03EB]=8'h65;
    mem['h03EC]=8'hBC; mem['h03ED]=8'hCD; mem['h03EE]=8'h98; mem['h03EF]=8'hD6;
    mem['h03F0]=8'h77; mem['h03F1]=8'h3E; mem['h03F2]=8'h98; mem['h03F3]=8'h52;
    mem['h03F4]=8'hC7; mem['h03F5]=8'h4F; mem['h03F6]=8'h80; mem['h03F7]=8'hDB;
    mem['h03F8]=8'h00; mem['h03F9]=8'hC9; mem['h03FA]=8'h01; mem['h03FB]=8'hFF;
    mem['h03FC]=8'h1C; mem['h03FD]=8'h00; mem['h03FE]=8'h00; mem['h03FF]=8'h14;
    mem['h0400]=8'h00; mem['h0401]=8'h14; mem['h0402]=8'h00; mem['h0403]=8'h00;
    mem['h0404]=8'h00; mem['h0405]=8'h00; mem['h0406]=8'h00; mem['h0407]=8'hC3;
    mem['h0408]=8'hCD; mem['h0409]=8'h06; mem['h040A]=8'hC3; mem['h040B]=8'h00;
    mem['h040C]=8'h00; mem['h040D]=8'hC3; mem['h040E]=8'h00; mem['h040F]=8'h00;
    mem['h0410]=8'hC3; mem['h0411]=8'h00; mem['h0412]=8'h00; mem['h0413]=8'hA2;
    mem['h0414]=8'h81; mem['h0415]=8'hFE; mem['h0416]=8'hFF; mem['h0417]=8'h3F;
    mem['h0418]=8'h81; mem['h0419]=8'h20; mem['h041A]=8'h45; mem['h041B]=8'h72;
    mem['h041C]=8'h72; mem['h041D]=8'h6F; mem['h041E]=8'h72; mem['h041F]=8'h00;
    mem['h0420]=8'h20; mem['h0421]=8'h69; mem['h0422]=8'h6E; mem['h0423]=8'h20;
    mem['h0424]=8'h00; mem['h0425]=8'h4F; mem['h0426]=8'h6B; mem['h0427]=8'h0D;
    mem['h0428]=8'h0A; mem['h0429]=8'h00; mem['h042A]=8'h00; mem['h042B]=8'h42;
    mem['h042C]=8'h72; mem['h042D]=8'h65; mem['h042E]=8'h61; mem['h042F]=8'h6B;
    mem['h0430]=8'h00; mem['h0431]=8'h21; mem['h0432]=8'h04; mem['h0433]=8'h00;
    mem['h0434]=8'h39; mem['h0435]=8'h7E; mem['h0436]=8'h23; mem['h0437]=8'hFE;
    mem['h0438]=8'h81; mem['h0439]=8'hC0; mem['h043A]=8'h4E; mem['h043B]=8'h23;
    mem['h043C]=8'h46; mem['h043D]=8'h23; mem['h043E]=8'hE5; mem['h043F]=8'h69;
    mem['h0440]=8'h60; mem['h0441]=8'h7A; mem['h0442]=8'hB3; mem['h0443]=8'hEB;
    mem['h0444]=8'hCA; mem['h0445]=8'h4B; mem['h0446]=8'h04; mem['h0447]=8'hEB;
    mem['h0448]=8'hCD; mem['h0449]=8'h50; mem['h044A]=8'h07; mem['h044B]=8'h01;
    mem['h044C]=8'h0D; mem['h044D]=8'h00; mem['h044E]=8'hE1; mem['h044F]=8'hC8;
    mem['h0450]=8'h09; mem['h0451]=8'hC3; mem['h0452]=8'h35; mem['h0453]=8'h04;
    mem['h0454]=8'hCD; mem['h0455]=8'h6E; mem['h0456]=8'h04; mem['h0457]=8'hC5;
    mem['h0458]=8'hE3; mem['h0459]=8'hC1; mem['h045A]=8'hCD; mem['h045B]=8'h50;
    mem['h045C]=8'h07; mem['h045D]=8'h7E; mem['h045E]=8'h02; mem['h045F]=8'hC8;
    mem['h0460]=8'h0B; mem['h0461]=8'h2B; mem['h0462]=8'hC3; mem['h0463]=8'h5A;
    mem['h0464]=8'h04; mem['h0465]=8'hE5; mem['h0466]=8'h2A; mem['h0467]=8'h1F;
    mem['h0468]=8'h81; mem['h0469]=8'h06; mem['h046A]=8'h00; mem['h046B]=8'h09;
    mem['h046C]=8'h09; mem['h046D]=8'h3E; mem['h046E]=8'hE5; mem['h046F]=8'h3E;
    mem['h0470]=8'hD0; mem['h0471]=8'h95; mem['h0472]=8'h6F; mem['h0473]=8'h3E;
    mem['h0474]=8'hFF; mem['h0475]=8'h9C; mem['h0476]=8'hDA; mem['h0477]=8'h7D;
    mem['h0478]=8'h04; mem['h0479]=8'h67; mem['h047A]=8'h39; mem['h047B]=8'hE1;
    mem['h047C]=8'hD8; mem['h047D]=8'h1E; mem['h047E]=8'h0C; mem['h047F]=8'hC3;
    mem['h0480]=8'h9C; mem['h0481]=8'h04; mem['h0482]=8'h2A; mem['h0483]=8'h0E;
    mem['h0484]=8'h81; mem['h0485]=8'h22; mem['h0486]=8'hA1; mem['h0487]=8'h80;
    mem['h0488]=8'h1E; mem['h0489]=8'h02; mem['h048A]=8'h01; mem['h048B]=8'h1E;
    mem['h048C]=8'h14; mem['h048D]=8'h01; mem['h048E]=8'h1E; mem['h048F]=8'h00;
    mem['h0490]=8'h01; mem['h0491]=8'h1E; mem['h0492]=8'h12; mem['h0493]=8'h01;
    mem['h0494]=8'h1E; mem['h0495]=8'h22; mem['h0496]=8'h01; mem['h0497]=8'h1E;
    mem['h0498]=8'h0A; mem['h0499]=8'h01; mem['h049A]=8'h1E; mem['h049B]=8'h18;
    mem['h049C]=8'hCD; mem['h049D]=8'hBA; mem['h049E]=8'h05; mem['h049F]=8'h32;
    mem['h04A0]=8'h8A; mem['h04A1]=8'h80; mem['h04A2]=8'hCD; mem['h04A3]=8'h7B;
    mem['h04A4]=8'h0B; mem['h04A5]=8'h21; mem['h04A6]=8'h8F; mem['h04A7]=8'h03;
    mem['h04A8]=8'h57; mem['h04A9]=8'h3E; mem['h04AA]=8'h3F; mem['h04AB]=8'hCD;
    mem['h04AC]=8'h61; mem['h04AD]=8'h07; mem['h04AE]=8'h19; mem['h04AF]=8'h7E;
    mem['h04B0]=8'hCD; mem['h04B1]=8'h61; mem['h04B2]=8'h07; mem['h04B3]=8'hCD;
    mem['h04B4]=8'hE0; mem['h04B5]=8'h08; mem['h04B6]=8'hCD; mem['h04B7]=8'h61;
    mem['h04B8]=8'h07; mem['h04B9]=8'h21; mem['h04BA]=8'h19; mem['h04BB]=8'h04;
    mem['h04BC]=8'hCD; mem['h04BD]=8'h26; mem['h04BE]=8'h12; mem['h04BF]=8'h2A;
    mem['h04C0]=8'hA1; mem['h04C1]=8'h80; mem['h04C2]=8'h11; mem['h04C3]=8'hFE;
    mem['h04C4]=8'hFF; mem['h04C5]=8'hCD; mem['h04C6]=8'h50; mem['h04C7]=8'h07;
    mem['h04C8]=8'hCA; mem['h04C9]=8'hE1; mem['h04CA]=8'h00; mem['h04CB]=8'h7C;
    mem['h04CC]=8'hA5; mem['h04CD]=8'h3C; mem['h04CE]=8'hC4; mem['h04CF]=8'hC1;
    mem['h04D0]=8'h18; mem['h04D1]=8'h3E; mem['h04D2]=8'hC1; mem['h04D3]=8'hAF;
    mem['h04D4]=8'h32; mem['h04D5]=8'h8A; mem['h04D6]=8'h80; mem['h04D7]=8'hCD;
    mem['h04D8]=8'h7B; mem['h04D9]=8'h0B; mem['h04DA]=8'h21; mem['h04DB]=8'h25;
    mem['h04DC]=8'h04; mem['h04DD]=8'hCD; mem['h04DE]=8'h26; mem['h04DF]=8'h12;
    mem['h04E0]=8'h21; mem['h04E1]=8'hFF; mem['h04E2]=8'hFF; mem['h04E3]=8'h22;
    mem['h04E4]=8'hA1; mem['h04E5]=8'h80; mem['h04E6]=8'hCD; mem['h04E7]=8'hCD;
    mem['h04E8]=8'h06; mem['h04E9]=8'hDA; mem['h04EA]=8'hE0; mem['h04EB]=8'h04;
    mem['h04EC]=8'hCD; mem['h04ED]=8'hE0; mem['h04EE]=8'h08; mem['h04EF]=8'h3C;
    mem['h04F0]=8'h3D; mem['h04F1]=8'hCA; mem['h04F2]=8'hE0; mem['h04F3]=8'h04;
    mem['h04F4]=8'hF5; mem['h04F5]=8'hCD; mem['h04F6]=8'hAC; mem['h04F7]=8'h09;
    mem['h04F8]=8'hD5; mem['h04F9]=8'hCD; mem['h04FA]=8'hE4; mem['h04FB]=8'h05;
    mem['h04FC]=8'h47; mem['h04FD]=8'hD1; mem['h04FE]=8'hF1; mem['h04FF]=8'hD2;
    mem['h0500]=8'hC0; mem['h0501]=8'h08; mem['h0502]=8'hD5; mem['h0503]=8'hC5;
    mem['h0504]=8'hAF; mem['h0505]=8'h32; mem['h0506]=8'h11; mem['h0507]=8'h81;
    mem['h0508]=8'hCD; mem['h0509]=8'hE0; mem['h050A]=8'h08; mem['h050B]=8'hB7;
    mem['h050C]=8'hF5; mem['h050D]=8'hCD; mem['h050E]=8'h74; mem['h050F]=8'h05;
    mem['h0510]=8'hDA; mem['h0511]=8'h19; mem['h0512]=8'h05; mem['h0513]=8'hF1;
    mem['h0514]=8'hF5; mem['h0515]=8'hCA; mem['h0516]=8'h4D; mem['h0517]=8'h0A;
    mem['h0518]=8'hB7; mem['h0519]=8'hC5; mem['h051A]=8'hD2; mem['h051B]=8'h30;
    mem['h051C]=8'h05; mem['h051D]=8'hEB; mem['h051E]=8'h2A; mem['h051F]=8'h1B;
    mem['h0520]=8'h81; mem['h0521]=8'h1A; mem['h0522]=8'h02; mem['h0523]=8'h03;
    mem['h0524]=8'h13; mem['h0525]=8'hCD; mem['h0526]=8'h50; mem['h0527]=8'h07;
    mem['h0528]=8'hC2; mem['h0529]=8'h21; mem['h052A]=8'h05; mem['h052B]=8'h60;
    mem['h052C]=8'h69; mem['h052D]=8'h22; mem['h052E]=8'h1B; mem['h052F]=8'h81;
    mem['h0530]=8'hD1; mem['h0531]=8'hF1; mem['h0532]=8'hCA; mem['h0533]=8'h57;
    mem['h0534]=8'h05; mem['h0535]=8'h2A; mem['h0536]=8'h1B; mem['h0537]=8'h81;
    mem['h0538]=8'hE3; mem['h0539]=8'hC1; mem['h053A]=8'h09; mem['h053B]=8'hE5;
    mem['h053C]=8'hCD; mem['h053D]=8'h54; mem['h053E]=8'h04; mem['h053F]=8'hE1;
    mem['h0540]=8'h22; mem['h0541]=8'h1B; mem['h0542]=8'h81; mem['h0543]=8'hEB;
    mem['h0544]=8'h74; mem['h0545]=8'hD1; mem['h0546]=8'h23; mem['h0547]=8'h23;
    mem['h0548]=8'h73; mem['h0549]=8'h23; mem['h054A]=8'h72; mem['h054B]=8'h23;
    mem['h054C]=8'h11; mem['h054D]=8'hA6; mem['h054E]=8'h80; mem['h054F]=8'h1A;
    mem['h0550]=8'h77; mem['h0551]=8'h23; mem['h0552]=8'h13; mem['h0553]=8'hB7;
    mem['h0554]=8'hC2; mem['h0555]=8'h4F; mem['h0556]=8'h05; mem['h0557]=8'hCD;
    mem['h0558]=8'hA0; mem['h0559]=8'h05; mem['h055A]=8'h23; mem['h055B]=8'hEB;
    mem['h055C]=8'h62; mem['h055D]=8'h6B; mem['h055E]=8'h7E; mem['h055F]=8'h23;
    mem['h0560]=8'hB6; mem['h0561]=8'hCA; mem['h0562]=8'hE0; mem['h0563]=8'h04;
    mem['h0564]=8'h23; mem['h0565]=8'h23; mem['h0566]=8'h23; mem['h0567]=8'hAF;
    mem['h0568]=8'hBE; mem['h0569]=8'h23; mem['h056A]=8'hC2; mem['h056B]=8'h68;
    mem['h056C]=8'h05; mem['h056D]=8'hEB; mem['h056E]=8'h73; mem['h056F]=8'h23;
    mem['h0570]=8'h72; mem['h0571]=8'hC3; mem['h0572]=8'h5C; mem['h0573]=8'h05;
    mem['h0574]=8'h2A; mem['h0575]=8'hA3; mem['h0576]=8'h80; mem['h0577]=8'h44;
    mem['h0578]=8'h4D; mem['h0579]=8'h7E; mem['h057A]=8'h23; mem['h057B]=8'hB6;
    mem['h057C]=8'h2B; mem['h057D]=8'hC8; mem['h057E]=8'h23; mem['h057F]=8'h23;
    mem['h0580]=8'h7E; mem['h0581]=8'h23; mem['h0582]=8'h66; mem['h0583]=8'h6F;
    mem['h0584]=8'hCD; mem['h0585]=8'h50; mem['h0586]=8'h07; mem['h0587]=8'h60;
    mem['h0588]=8'h69; mem['h0589]=8'h7E; mem['h058A]=8'h23; mem['h058B]=8'h66;
    mem['h058C]=8'h6F; mem['h058D]=8'h3F; mem['h058E]=8'hC8; mem['h058F]=8'h3F;
    mem['h0590]=8'hD0; mem['h0591]=8'hC3; mem['h0592]=8'h77; mem['h0593]=8'h05;
    mem['h0594]=8'hC0; mem['h0595]=8'h2A; mem['h0596]=8'hA3; mem['h0597]=8'h80;
    mem['h0598]=8'hAF; mem['h0599]=8'h77; mem['h059A]=8'h23; mem['h059B]=8'h77;
    mem['h059C]=8'h23; mem['h059D]=8'h22; mem['h059E]=8'h1B; mem['h059F]=8'h81;
    mem['h05A0]=8'h2A; mem['h05A1]=8'hA3; mem['h05A2]=8'h80; mem['h05A3]=8'h2B;
    mem['h05A4]=8'h22; mem['h05A5]=8'h13; mem['h05A6]=8'h81; mem['h05A7]=8'h2A;
    mem['h05A8]=8'hF4; mem['h05A9]=8'h80; mem['h05AA]=8'h22; mem['h05AB]=8'h08;
    mem['h05AC]=8'h81; mem['h05AD]=8'hAF; mem['h05AE]=8'hCD; mem['h05AF]=8'hF0;
    mem['h05B0]=8'h08; mem['h05B1]=8'h2A; mem['h05B2]=8'h1B; mem['h05B3]=8'h81;
    mem['h05B4]=8'h22; mem['h05B5]=8'h1D; mem['h05B6]=8'h81; mem['h05B7]=8'h22;
    mem['h05B8]=8'h1F; mem['h05B9]=8'h81; mem['h05BA]=8'hC1; mem['h05BB]=8'h2A;
    mem['h05BC]=8'h9F; mem['h05BD]=8'h80; mem['h05BE]=8'hF9; mem['h05BF]=8'h21;
    mem['h05C0]=8'hF8; mem['h05C1]=8'h80; mem['h05C2]=8'h22; mem['h05C3]=8'hF6;
    mem['h05C4]=8'h80; mem['h05C5]=8'hAF; mem['h05C6]=8'h6F; mem['h05C7]=8'h67;
    mem['h05C8]=8'h22; mem['h05C9]=8'h19; mem['h05CA]=8'h81; mem['h05CB]=8'h32;
    mem['h05CC]=8'h10; mem['h05CD]=8'h81; mem['h05CE]=8'h22; mem['h05CF]=8'h23;
    mem['h05D0]=8'h81; mem['h05D1]=8'hE5; mem['h05D2]=8'hC5; mem['h05D3]=8'h2A;
    mem['h05D4]=8'h13; mem['h05D5]=8'h81; mem['h05D6]=8'hC9; mem['h05D7]=8'h3E;
    mem['h05D8]=8'h3F; mem['h05D9]=8'hCD; mem['h05DA]=8'h61; mem['h05DB]=8'h07;
    mem['h05DC]=8'h3E; mem['h05DD]=8'h20; mem['h05DE]=8'hCD; mem['h05DF]=8'h61;
    mem['h05E0]=8'h07; mem['h05E1]=8'hC3; mem['h05E2]=8'h93; mem['h05E3]=8'h80;
    mem['h05E4]=8'hAF; mem['h05E5]=8'h32; mem['h05E6]=8'hF3; mem['h05E7]=8'h80;
    mem['h05E8]=8'h0E; mem['h05E9]=8'h05; mem['h05EA]=8'h11; mem['h05EB]=8'hA6;
    mem['h05EC]=8'h80; mem['h05ED]=8'h7E; mem['h05EE]=8'hFE; mem['h05EF]=8'h20;
    mem['h05F0]=8'hCA; mem['h05F1]=8'h6C; mem['h05F2]=8'h06; mem['h05F3]=8'h47;
    mem['h05F4]=8'hFE; mem['h05F5]=8'h22; mem['h05F6]=8'hCA; mem['h05F7]=8'h8C;
    mem['h05F8]=8'h06; mem['h05F9]=8'hB7; mem['h05FA]=8'hCA; mem['h05FB]=8'h93;
    mem['h05FC]=8'h06; mem['h05FD]=8'h3A; mem['h05FE]=8'hF3; mem['h05FF]=8'h80;
    mem['h0600]=8'hB7; mem['h0601]=8'h7E; mem['h0602]=8'hC2; mem['h0603]=8'h6C;
    mem['h0604]=8'h06; mem['h0605]=8'hFE; mem['h0606]=8'h3F; mem['h0607]=8'h3E;
    mem['h0608]=8'h9E; mem['h0609]=8'hCA; mem['h060A]=8'h6C; mem['h060B]=8'h06;
    mem['h060C]=8'h7E; mem['h060D]=8'hFE; mem['h060E]=8'h30; mem['h060F]=8'hDA;
    mem['h0610]=8'h17; mem['h0611]=8'h06; mem['h0612]=8'hFE; mem['h0613]=8'h3C;
    mem['h0614]=8'hDA; mem['h0615]=8'h6C; mem['h0616]=8'h06; mem['h0617]=8'hD5;
    mem['h0618]=8'h11; mem['h0619]=8'h10; mem['h061A]=8'h02; mem['h061B]=8'hC5;
    mem['h061C]=8'h01; mem['h061D]=8'h68; mem['h061E]=8'h06; mem['h061F]=8'hC5;
    mem['h0620]=8'h06; mem['h0621]=8'h7F; mem['h0622]=8'h7E; mem['h0623]=8'hFE;
    mem['h0624]=8'h61; mem['h0625]=8'hDA; mem['h0626]=8'h30; mem['h0627]=8'h06;
    mem['h0628]=8'hFE; mem['h0629]=8'h7B; mem['h062A]=8'hD2; mem['h062B]=8'h30;
    mem['h062C]=8'h06; mem['h062D]=8'hE6; mem['h062E]=8'h5F; mem['h062F]=8'h77;
    mem['h0630]=8'h4E; mem['h0631]=8'hEB; mem['h0632]=8'h23; mem['h0633]=8'hB6;
    mem['h0634]=8'hF2; mem['h0635]=8'h32; mem['h0636]=8'h06; mem['h0637]=8'h04;
    mem['h0638]=8'h7E; mem['h0639]=8'hE6; mem['h063A]=8'h7F; mem['h063B]=8'hC8;
    mem['h063C]=8'hB9; mem['h063D]=8'hC2; mem['h063E]=8'h32; mem['h063F]=8'h06;
    mem['h0640]=8'hEB; mem['h0641]=8'hE5; mem['h0642]=8'h13; mem['h0643]=8'h1A;
    mem['h0644]=8'hB7; mem['h0645]=8'hFA; mem['h0646]=8'h64; mem['h0647]=8'h06;
    mem['h0648]=8'h4F; mem['h0649]=8'h78; mem['h064A]=8'hFE; mem['h064B]=8'h88;
    mem['h064C]=8'hC2; mem['h064D]=8'h53; mem['h064E]=8'h06; mem['h064F]=8'hCD;
    mem['h0650]=8'hE0; mem['h0651]=8'h08; mem['h0652]=8'h2B; mem['h0653]=8'h23;
    mem['h0654]=8'h7E; mem['h0655]=8'hFE; mem['h0656]=8'h61; mem['h0657]=8'hDA;
    mem['h0658]=8'h5C; mem['h0659]=8'h06; mem['h065A]=8'hE6; mem['h065B]=8'h5F;
    mem['h065C]=8'hB9; mem['h065D]=8'hCA; mem['h065E]=8'h42; mem['h065F]=8'h06;
    mem['h0660]=8'hE1; mem['h0661]=8'hC3; mem['h0662]=8'h30; mem['h0663]=8'h06;
    mem['h0664]=8'h48; mem['h0665]=8'hF1; mem['h0666]=8'hEB; mem['h0667]=8'hC9;
    mem['h0668]=8'hEB; mem['h0669]=8'h79; mem['h066A]=8'hC1; mem['h066B]=8'hD1;
    mem['h066C]=8'h23; mem['h066D]=8'h12; mem['h066E]=8'h13; mem['h066F]=8'h0C;
    mem['h0670]=8'hD6; mem['h0671]=8'h3A; mem['h0672]=8'hCA; mem['h0673]=8'h7A;
    mem['h0674]=8'h06; mem['h0675]=8'hFE; mem['h0676]=8'h49; mem['h0677]=8'hC2;
    mem['h0678]=8'h7D; mem['h0679]=8'h06; mem['h067A]=8'h32; mem['h067B]=8'hF3;
    mem['h067C]=8'h80; mem['h067D]=8'hD6; mem['h067E]=8'h54; mem['h067F]=8'hC2;
    mem['h0680]=8'hED; mem['h0681]=8'h05; mem['h0682]=8'h47; mem['h0683]=8'h7E;
    mem['h0684]=8'hB7; mem['h0685]=8'hCA; mem['h0686]=8'h93; mem['h0687]=8'h06;
    mem['h0688]=8'hB8; mem['h0689]=8'hCA; mem['h068A]=8'h6C; mem['h068B]=8'h06;
    mem['h068C]=8'h23; mem['h068D]=8'h12; mem['h068E]=8'h0C; mem['h068F]=8'h13;
    mem['h0690]=8'hC3; mem['h0691]=8'h83; mem['h0692]=8'h06; mem['h0693]=8'h21;
    mem['h0694]=8'hA5; mem['h0695]=8'h80; mem['h0696]=8'h12; mem['h0697]=8'h13;
    mem['h0698]=8'h12; mem['h0699]=8'h13; mem['h069A]=8'h12; mem['h069B]=8'hC9;
    mem['h069C]=8'h3A; mem['h069D]=8'h89; mem['h069E]=8'h80; mem['h069F]=8'hB7;
    mem['h06A0]=8'h3E; mem['h06A1]=8'h00; mem['h06A2]=8'h32; mem['h06A3]=8'h89;
    mem['h06A4]=8'h80; mem['h06A5]=8'hC2; mem['h06A6]=8'hB0; mem['h06A7]=8'h06;
    mem['h06A8]=8'h05; mem['h06A9]=8'hCA; mem['h06AA]=8'hCD; mem['h06AB]=8'h06;
    mem['h06AC]=8'hCD; mem['h06AD]=8'h61; mem['h06AE]=8'h07; mem['h06AF]=8'h3E;
    mem['h06B0]=8'h05; mem['h06B1]=8'h2B; mem['h06B2]=8'hCA; mem['h06B3]=8'hC4;
    mem['h06B4]=8'h06; mem['h06B5]=8'h7E; mem['h06B6]=8'hCD; mem['h06B7]=8'h61;
    mem['h06B8]=8'h07; mem['h06B9]=8'hC3; mem['h06BA]=8'hD6; mem['h06BB]=8'h06;
    mem['h06BC]=8'h05; mem['h06BD]=8'h2B; mem['h06BE]=8'hCD; mem['h06BF]=8'h61;
    mem['h06C0]=8'h07; mem['h06C1]=8'hC2; mem['h06C2]=8'hD6; mem['h06C3]=8'h06;
    mem['h06C4]=8'hCD; mem['h06C5]=8'h61; mem['h06C6]=8'h07; mem['h06C7]=8'hCD;
    mem['h06C8]=8'h88; mem['h06C9]=8'h0B; mem['h06CA]=8'hC3; mem['h06CB]=8'hCD;
    mem['h06CC]=8'h06; mem['h06CD]=8'h21; mem['h06CE]=8'hA6; mem['h06CF]=8'h80;
    mem['h06D0]=8'h06; mem['h06D1]=8'h01; mem['h06D2]=8'hAF; mem['h06D3]=8'h32;
    mem['h06D4]=8'h89; mem['h06D5]=8'h80; mem['h06D6]=8'hCD; mem['h06D7]=8'h8B;
    mem['h06D8]=8'h07; mem['h06D9]=8'h4F; mem['h06DA]=8'hFE; mem['h06DB]=8'h7F;
    mem['h06DC]=8'hCA; mem['h06DD]=8'h9C; mem['h06DE]=8'h06; mem['h06DF]=8'h3A;
    mem['h06E0]=8'h89; mem['h06E1]=8'h80; mem['h06E2]=8'hB7; mem['h06E3]=8'hCA;
    mem['h06E4]=8'hEF; mem['h06E5]=8'h06; mem['h06E6]=8'h3E; mem['h06E7]=8'h00;
    mem['h06E8]=8'hCD; mem['h06E9]=8'h61; mem['h06EA]=8'h07; mem['h06EB]=8'hAF;
    mem['h06EC]=8'h32; mem['h06ED]=8'h89; mem['h06EE]=8'h80; mem['h06EF]=8'h79;
    mem['h06F0]=8'hFE; mem['h06F1]=8'h07; mem['h06F2]=8'hCA; mem['h06F3]=8'h33;
    mem['h06F4]=8'h07; mem['h06F5]=8'hFE; mem['h06F6]=8'h03; mem['h06F7]=8'hCC;
    mem['h06F8]=8'h88; mem['h06F9]=8'h0B; mem['h06FA]=8'h37; mem['h06FB]=8'hC8;
    mem['h06FC]=8'hFE; mem['h06FD]=8'h0D; mem['h06FE]=8'hCA; mem['h06FF]=8'h83;
    mem['h0700]=8'h0B; mem['h0701]=8'hFE; mem['h0702]=8'h15; mem['h0703]=8'hCA;
    mem['h0704]=8'hC7; mem['h0705]=8'h06; mem['h0706]=8'hFE; mem['h0707]=8'h40;
    mem['h0708]=8'hCA; mem['h0709]=8'hC4; mem['h070A]=8'h06; mem['h070B]=8'hFE;
    mem['h070C]=8'h5F; mem['h070D]=8'hCA; mem['h070E]=8'hBC; mem['h070F]=8'h06;
    mem['h0710]=8'hFE; mem['h0711]=8'h08; mem['h0712]=8'hCA; mem['h0713]=8'hBC;
    mem['h0714]=8'h06; mem['h0715]=8'hFE; mem['h0716]=8'h12; mem['h0717]=8'hC2;
    mem['h0718]=8'h2E; mem['h0719]=8'h07; mem['h071A]=8'hC5; mem['h071B]=8'hD5;
    mem['h071C]=8'hE5; mem['h071D]=8'h36; mem['h071E]=8'h00; mem['h071F]=8'hCD;
    mem['h0720]=8'h32; mem['h0721]=8'h1D; mem['h0722]=8'h21; mem['h0723]=8'hA6;
    mem['h0724]=8'h80; mem['h0725]=8'hCD; mem['h0726]=8'h26; mem['h0727]=8'h12;
    mem['h0728]=8'hE1; mem['h0729]=8'hD1; mem['h072A]=8'hC1; mem['h072B]=8'hC3;
    mem['h072C]=8'hD6; mem['h072D]=8'h06; mem['h072E]=8'hFE; mem['h072F]=8'h20;
    mem['h0730]=8'hDA; mem['h0731]=8'hD6; mem['h0732]=8'h06; mem['h0733]=8'h78;
    mem['h0734]=8'hFE; mem['h0735]=8'h49; mem['h0736]=8'h3E; mem['h0737]=8'h07;
    mem['h0738]=8'hD2; mem['h0739]=8'h48; mem['h073A]=8'h07; mem['h073B]=8'h79;
    mem['h073C]=8'h71; mem['h073D]=8'h32; mem['h073E]=8'h11; mem['h073F]=8'h81;
    mem['h0740]=8'h23; mem['h0741]=8'h04; mem['h0742]=8'hCD; mem['h0743]=8'h61;
    mem['h0744]=8'h07; mem['h0745]=8'hC3; mem['h0746]=8'hD6; mem['h0747]=8'h06;
    mem['h0748]=8'hCD; mem['h0749]=8'h61; mem['h074A]=8'h07; mem['h074B]=8'h3E;
    mem['h074C]=8'h08; mem['h074D]=8'hC3; mem['h074E]=8'h42; mem['h074F]=8'h07;
    mem['h0750]=8'h7C; mem['h0751]=8'h92; mem['h0752]=8'hC0; mem['h0753]=8'h7D;
    mem['h0754]=8'h93; mem['h0755]=8'hC9; mem['h0756]=8'h7E; mem['h0757]=8'hE3;
    mem['h0758]=8'hBE; mem['h0759]=8'h23; mem['h075A]=8'hE3; mem['h075B]=8'hCA;
    mem['h075C]=8'hE0; mem['h075D]=8'h08; mem['h075E]=8'hC3; mem['h075F]=8'h88;
    mem['h0760]=8'h04; mem['h0761]=8'hF5; mem['h0762]=8'h3A; mem['h0763]=8'h8A;
    mem['h0764]=8'h80; mem['h0765]=8'hB7; mem['h0766]=8'hC2; mem['h0767]=8'h5B;
    mem['h0768]=8'h12; mem['h0769]=8'hF1; mem['h076A]=8'hC5; mem['h076B]=8'hF5;
    mem['h076C]=8'hFE; mem['h076D]=8'h20; mem['h076E]=8'hDA; mem['h076F]=8'h85;
    mem['h0770]=8'h07; mem['h0771]=8'h3A; mem['h0772]=8'h87; mem['h0773]=8'h80;
    mem['h0774]=8'h47; mem['h0775]=8'h3A; mem['h0776]=8'hF0; mem['h0777]=8'h80;
    mem['h0778]=8'h04; mem['h0779]=8'hCA; mem['h077A]=8'h81; mem['h077B]=8'h07;
    mem['h077C]=8'h05; mem['h077D]=8'hB8; mem['h077E]=8'hCC; mem['h077F]=8'h88;
    mem['h0780]=8'h0B; mem['h0781]=8'h3C; mem['h0782]=8'h32; mem['h0783]=8'hF0;
    mem['h0784]=8'h80; mem['h0785]=8'hF1; mem['h0786]=8'hC1; mem['h0787]=8'hCD;
    mem['h0788]=8'h1D; mem['h0789]=8'h1D; mem['h078A]=8'hC9; mem['h078B]=8'hCD;
    mem['h078C]=8'hE5; mem['h078D]=8'h1B; mem['h078E]=8'hE6; mem['h078F]=8'h7F;
    mem['h0790]=8'hFE; mem['h0791]=8'h0F; mem['h0792]=8'hC0; mem['h0793]=8'h3A;
    mem['h0794]=8'h8A; mem['h0795]=8'h80; mem['h0796]=8'h2F; mem['h0797]=8'h32;
    mem['h0798]=8'h8A; mem['h0799]=8'h80; mem['h079A]=8'hAF; mem['h079B]=8'hC9;
    mem['h079C]=8'hCD; mem['h079D]=8'hAC; mem['h079E]=8'h09; mem['h079F]=8'hC0;
    mem['h07A0]=8'hC1; mem['h07A1]=8'hCD; mem['h07A2]=8'h74; mem['h07A3]=8'h05;
    mem['h07A4]=8'hC5; mem['h07A5]=8'hCD; mem['h07A6]=8'hF2; mem['h07A7]=8'h07;
    mem['h07A8]=8'hE1; mem['h07A9]=8'h4E; mem['h07AA]=8'h23; mem['h07AB]=8'h46;
    mem['h07AC]=8'h23; mem['h07AD]=8'h78; mem['h07AE]=8'hB1; mem['h07AF]=8'hCA;
    mem['h07B0]=8'hD3; mem['h07B1]=8'h04; mem['h07B2]=8'hCD; mem['h07B3]=8'hFB;
    mem['h07B4]=8'h07; mem['h07B5]=8'hCD; mem['h07B6]=8'h0B; mem['h07B7]=8'h09;
    mem['h07B8]=8'hC5; mem['h07B9]=8'hCD; mem['h07BA]=8'h88; mem['h07BB]=8'h0B;
    mem['h07BC]=8'h5E; mem['h07BD]=8'h23; mem['h07BE]=8'h56; mem['h07BF]=8'h23;
    mem['h07C0]=8'hE5; mem['h07C1]=8'hEB; mem['h07C2]=8'hCD; mem['h07C3]=8'hC9;
    mem['h07C4]=8'h18; mem['h07C5]=8'h3E; mem['h07C6]=8'h20; mem['h07C7]=8'hE1;
    mem['h07C8]=8'hCD; mem['h07C9]=8'h61; mem['h07CA]=8'h07; mem['h07CB]=8'h7E;
    mem['h07CC]=8'hB7; mem['h07CD]=8'h23; mem['h07CE]=8'hCA; mem['h07CF]=8'hA8;
    mem['h07D0]=8'h07; mem['h07D1]=8'hF2; mem['h07D2]=8'hC8; mem['h07D3]=8'h07;
    mem['h07D4]=8'hD6; mem['h07D5]=8'h7F; mem['h07D6]=8'h4F; mem['h07D7]=8'h11;
    mem['h07D8]=8'h11; mem['h07D9]=8'h02; mem['h07DA]=8'h1A; mem['h07DB]=8'h13;
    mem['h07DC]=8'hB7; mem['h07DD]=8'hF2; mem['h07DE]=8'hDA; mem['h07DF]=8'h07;
    mem['h07E0]=8'h0D; mem['h07E1]=8'hC2; mem['h07E2]=8'hDA; mem['h07E3]=8'h07;
    mem['h07E4]=8'hE6; mem['h07E5]=8'h7F; mem['h07E6]=8'hCD; mem['h07E7]=8'h61;
    mem['h07E8]=8'h07; mem['h07E9]=8'h1A; mem['h07EA]=8'h13; mem['h07EB]=8'hB7;
    mem['h07EC]=8'hF2; mem['h07ED]=8'hE4; mem['h07EE]=8'h07; mem['h07EF]=8'hC3;
    mem['h07F0]=8'hCB; mem['h07F1]=8'h07; mem['h07F2]=8'hE5; mem['h07F3]=8'h2A;
    mem['h07F4]=8'h8D; mem['h07F5]=8'h80; mem['h07F6]=8'h22; mem['h07F7]=8'h8B;
    mem['h07F8]=8'h80; mem['h07F9]=8'hE1; mem['h07FA]=8'hC9; mem['h07FB]=8'hE5;
    mem['h07FC]=8'hD5; mem['h07FD]=8'h2A; mem['h07FE]=8'h8B; mem['h07FF]=8'h80;
    mem['h0800]=8'h11; mem['h0801]=8'hFF; mem['h0802]=8'hFF; mem['h0803]=8'hED;
    mem['h0804]=8'h5A; mem['h0805]=8'h22; mem['h0806]=8'h8B; mem['h0807]=8'h80;
    mem['h0808]=8'hD1; mem['h0809]=8'hE1; mem['h080A]=8'hF0; mem['h080B]=8'hE5;
    mem['h080C]=8'h2A; mem['h080D]=8'h8D; mem['h080E]=8'h80; mem['h080F]=8'h22;
    mem['h0810]=8'h8B; mem['h0811]=8'h80; mem['h0812]=8'hCD; mem['h0813]=8'hE5;
    mem['h0814]=8'h1B; mem['h0815]=8'hFE; mem['h0816]=8'h03; mem['h0817]=8'hCA;
    mem['h0818]=8'h1E; mem['h0819]=8'h08; mem['h081A]=8'hE1; mem['h081B]=8'hC3;
    mem['h081C]=8'hFB; mem['h081D]=8'h07; mem['h081E]=8'h2A; mem['h081F]=8'h8D;
    mem['h0820]=8'h80; mem['h0821]=8'h22; mem['h0822]=8'h8B; mem['h0823]=8'h80;
    mem['h0824]=8'hC3; mem['h0825]=8'h52; mem['h0826]=8'h01; mem['h0827]=8'h3E;
    mem['h0828]=8'h64; mem['h0829]=8'h32; mem['h082A]=8'h10; mem['h082B]=8'h81;
    mem['h082C]=8'hCD; mem['h082D]=8'h8E; mem['h082E]=8'h0A; mem['h082F]=8'hC1;
    mem['h0830]=8'hE5; mem['h0831]=8'hCD; mem['h0832]=8'h77; mem['h0833]=8'h0A;
    mem['h0834]=8'h22; mem['h0835]=8'h0C; mem['h0836]=8'h81; mem['h0837]=8'h21;
    mem['h0838]=8'h02; mem['h0839]=8'h00; mem['h083A]=8'h39; mem['h083B]=8'hCD;
    mem['h083C]=8'h35; mem['h083D]=8'h04; mem['h083E]=8'hD1; mem['h083F]=8'hC2;
    mem['h0840]=8'h57; mem['h0841]=8'h08; mem['h0842]=8'h09; mem['h0843]=8'hD5;
    mem['h0844]=8'h2B; mem['h0845]=8'h56; mem['h0846]=8'h2B; mem['h0847]=8'h5E;
    mem['h0848]=8'h23; mem['h0849]=8'h23; mem['h084A]=8'hE5; mem['h084B]=8'h2A;
    mem['h084C]=8'h0C; mem['h084D]=8'h81; mem['h084E]=8'hCD; mem['h084F]=8'h50;
    mem['h0850]=8'h07; mem['h0851]=8'hE1; mem['h0852]=8'hC2; mem['h0853]=8'h3B;
    mem['h0854]=8'h08; mem['h0855]=8'hD1; mem['h0856]=8'hF9; mem['h0857]=8'hEB;
    mem['h0858]=8'h0E; mem['h0859]=8'h08; mem['h085A]=8'hCD; mem['h085B]=8'h65;
    mem['h085C]=8'h04; mem['h085D]=8'hE5; mem['h085E]=8'h2A; mem['h085F]=8'h0C;
    mem['h0860]=8'h81; mem['h0861]=8'hE3; mem['h0862]=8'hE5; mem['h0863]=8'h2A;
    mem['h0864]=8'hA1; mem['h0865]=8'h80; mem['h0866]=8'hE3; mem['h0867]=8'hCD;
    mem['h0868]=8'h50; mem['h0869]=8'h0D; mem['h086A]=8'hCD; mem['h086B]=8'h56;
    mem['h086C]=8'h07; mem['h086D]=8'hA6; mem['h086E]=8'hCD; mem['h086F]=8'h4D;
    mem['h0870]=8'h0D; mem['h0871]=8'hE5; mem['h0872]=8'hCD; mem['h0873]=8'h7B;
    mem['h0874]=8'h17; mem['h0875]=8'hE1; mem['h0876]=8'hC5; mem['h0877]=8'hD5;
    mem['h0878]=8'h01; mem['h0879]=8'h00; mem['h087A]=8'h81; mem['h087B]=8'h51;
    mem['h087C]=8'h5A; mem['h087D]=8'h7E; mem['h087E]=8'hFE; mem['h087F]=8'hAB;
    mem['h0880]=8'h3E; mem['h0881]=8'h01; mem['h0882]=8'hC2; mem['h0883]=8'h93;
    mem['h0884]=8'h08; mem['h0885]=8'hCD; mem['h0886]=8'hE0; mem['h0887]=8'h08;
    mem['h0888]=8'hCD; mem['h0889]=8'h4D; mem['h088A]=8'h0D; mem['h088B]=8'hE5;
    mem['h088C]=8'hCD; mem['h088D]=8'h7B; mem['h088E]=8'h17; mem['h088F]=8'hCD;
    mem['h0890]=8'h2F; mem['h0891]=8'h17; mem['h0892]=8'hE1; mem['h0893]=8'hC5;
    mem['h0894]=8'hD5; mem['h0895]=8'hF5; mem['h0896]=8'h33; mem['h0897]=8'hE5;
    mem['h0898]=8'h2A; mem['h0899]=8'h13; mem['h089A]=8'h81; mem['h089B]=8'hE3;
    mem['h089C]=8'h06; mem['h089D]=8'h81; mem['h089E]=8'hC5; mem['h089F]=8'h33;
    mem['h08A0]=8'hCD; mem['h08A1]=8'h0B; mem['h08A2]=8'h09; mem['h08A3]=8'h22;
    mem['h08A4]=8'h13; mem['h08A5]=8'h81; mem['h08A6]=8'h7E; mem['h08A7]=8'hFE;
    mem['h08A8]=8'h3A; mem['h08A9]=8'hCA; mem['h08AA]=8'hC0; mem['h08AB]=8'h08;
    mem['h08AC]=8'hB7; mem['h08AD]=8'hC2; mem['h08AE]=8'h88; mem['h08AF]=8'h04;
    mem['h08B0]=8'h23; mem['h08B1]=8'h7E; mem['h08B2]=8'h23; mem['h08B3]=8'hB6;
    mem['h08B4]=8'hCA; mem['h08B5]=8'h32; mem['h08B6]=8'h09; mem['h08B7]=8'h23;
    mem['h08B8]=8'h5E; mem['h08B9]=8'h23; mem['h08BA]=8'h56; mem['h08BB]=8'hEB;
    mem['h08BC]=8'h22; mem['h08BD]=8'hA1; mem['h08BE]=8'h80; mem['h08BF]=8'hEB;
    mem['h08C0]=8'hCD; mem['h08C1]=8'hE0; mem['h08C2]=8'h08; mem['h08C3]=8'h11;
    mem['h08C4]=8'hA0; mem['h08C5]=8'h08; mem['h08C6]=8'hD5; mem['h08C7]=8'hC8;
    mem['h08C8]=8'hD6; mem['h08C9]=8'h80; mem['h08CA]=8'hDA; mem['h08CB]=8'h8E;
    mem['h08CC]=8'h0A; mem['h08CD]=8'hFE; mem['h08CE]=8'h25; mem['h08CF]=8'hD2;
    mem['h08D0]=8'h88; mem['h08D1]=8'h04; mem['h08D2]=8'h07; mem['h08D3]=8'h4F;
    mem['h08D4]=8'h06; mem['h08D5]=8'h00; mem['h08D6]=8'hEB; mem['h08D7]=8'h21;
    mem['h08D8]=8'h30; mem['h08D9]=8'h03; mem['h08DA]=8'h09; mem['h08DB]=8'h4E;
    mem['h08DC]=8'h23; mem['h08DD]=8'h46; mem['h08DE]=8'hC5; mem['h08DF]=8'hEB;
    mem['h08E0]=8'h23; mem['h08E1]=8'h7E; mem['h08E2]=8'hFE; mem['h08E3]=8'h3A;
    mem['h08E4]=8'hD0; mem['h08E5]=8'hFE; mem['h08E6]=8'h20; mem['h08E7]=8'hCA;
    mem['h08E8]=8'hE0; mem['h08E9]=8'h08; mem['h08EA]=8'hFE; mem['h08EB]=8'h30;
    mem['h08EC]=8'h3F; mem['h08ED]=8'h3C; mem['h08EE]=8'h3D; mem['h08EF]=8'hC9;
    mem['h08F0]=8'hEB; mem['h08F1]=8'h2A; mem['h08F2]=8'hA3; mem['h08F3]=8'h80;
    mem['h08F4]=8'hCA; mem['h08F5]=8'h05; mem['h08F6]=8'h09; mem['h08F7]=8'hEB;
    mem['h08F8]=8'hCD; mem['h08F9]=8'hAC; mem['h08FA]=8'h09; mem['h08FB]=8'hE5;
    mem['h08FC]=8'hCD; mem['h08FD]=8'h74; mem['h08FE]=8'h05; mem['h08FF]=8'h60;
    mem['h0900]=8'h69; mem['h0901]=8'hD1; mem['h0902]=8'hD2; mem['h0903]=8'h4D;
    mem['h0904]=8'h0A; mem['h0905]=8'h2B; mem['h0906]=8'h22; mem['h0907]=8'h21;
    mem['h0908]=8'h81; mem['h0909]=8'hEB; mem['h090A]=8'hC9; mem['h090B]=8'hDF;
    mem['h090C]=8'hC8; mem['h090D]=8'hD7; mem['h090E]=8'hFE; mem['h090F]=8'h1B;
    mem['h0910]=8'h28; mem['h0911]=8'h11; mem['h0912]=8'hFE; mem['h0913]=8'h03;
    mem['h0914]=8'h28; mem['h0915]=8'h0D; mem['h0916]=8'hFE; mem['h0917]=8'h13;
    mem['h0918]=8'hC0; mem['h0919]=8'hD7; mem['h091A]=8'hFE; mem['h091B]=8'h11;
    mem['h091C]=8'hC8; mem['h091D]=8'hFE; mem['h091E]=8'h03; mem['h091F]=8'h28;
    mem['h0920]=8'h07; mem['h0921]=8'h18; mem['h0922]=8'hF6; mem['h0923]=8'h3E;
    mem['h0924]=8'hFF; mem['h0925]=8'h32; mem['h0926]=8'h92; mem['h0927]=8'h80;
    mem['h0928]=8'hC0; mem['h0929]=8'hF6; mem['h092A]=8'hC0; mem['h092B]=8'h22;
    mem['h092C]=8'h13; mem['h092D]=8'h81; mem['h092E]=8'h21; mem['h092F]=8'hF6;
    mem['h0930]=8'hFF; mem['h0931]=8'hC1; mem['h0932]=8'h2A; mem['h0933]=8'hA1;
    mem['h0934]=8'h80; mem['h0935]=8'hF5; mem['h0936]=8'h7D; mem['h0937]=8'hA4;
    mem['h0938]=8'h3C; mem['h0939]=8'hCA; mem['h093A]=8'h45; mem['h093B]=8'h09;
    mem['h093C]=8'h22; mem['h093D]=8'h17; mem['h093E]=8'h81; mem['h093F]=8'h2A;
    mem['h0940]=8'h13; mem['h0941]=8'h81; mem['h0942]=8'h22; mem['h0943]=8'h19;
    mem['h0944]=8'h81; mem['h0945]=8'hAF; mem['h0946]=8'h32; mem['h0947]=8'h8A;
    mem['h0948]=8'h80; mem['h0949]=8'hCD; mem['h094A]=8'h7B; mem['h094B]=8'h0B;
    mem['h094C]=8'hF1; mem['h094D]=8'h21; mem['h094E]=8'h2B; mem['h094F]=8'h04;
    mem['h0950]=8'hC2; mem['h0951]=8'hBC; mem['h0952]=8'h04; mem['h0953]=8'hC3;
    mem['h0954]=8'hD3; mem['h0955]=8'h04; mem['h0956]=8'h2A; mem['h0957]=8'h19;
    mem['h0958]=8'h81; mem['h0959]=8'h7C; mem['h095A]=8'hB5; mem['h095B]=8'h1E;
    mem['h095C]=8'h20; mem['h095D]=8'hCA; mem['h095E]=8'h9C; mem['h095F]=8'h04;
    mem['h0960]=8'hEB; mem['h0961]=8'h2A; mem['h0962]=8'h17; mem['h0963]=8'h81;
    mem['h0964]=8'h22; mem['h0965]=8'hA1; mem['h0966]=8'h80; mem['h0967]=8'hEB;
    mem['h0968]=8'hC9; mem['h0969]=8'hCD; mem['h096A]=8'hAE; mem['h096B]=8'h14;
    mem['h096C]=8'hC0; mem['h096D]=8'h32; mem['h096E]=8'h86; mem['h096F]=8'h80;
    mem['h0970]=8'hC9; mem['h0971]=8'hE5; mem['h0972]=8'h2A; mem['h0973]=8'h8F;
    mem['h0974]=8'h80; mem['h0975]=8'h06; mem['h0976]=8'h00; mem['h0977]=8'h4F;
    mem['h0978]=8'h09; mem['h0979]=8'h22; mem['h097A]=8'h8F; mem['h097B]=8'h80;
    mem['h097C]=8'hE1; mem['h097D]=8'hC9; mem['h097E]=8'h7E; mem['h097F]=8'hFE;
    mem['h0980]=8'h41; mem['h0981]=8'hD8; mem['h0982]=8'hFE; mem['h0983]=8'h5B;
    mem['h0984]=8'h3F; mem['h0985]=8'hC9; mem['h0986]=8'hCD; mem['h0987]=8'hE0;
    mem['h0988]=8'h08; mem['h0989]=8'hCD; mem['h098A]=8'h4D; mem['h098B]=8'h0D;
    mem['h098C]=8'hCD; mem['h098D]=8'h2F; mem['h098E]=8'h17; mem['h098F]=8'hFA;
    mem['h0990]=8'hA7; mem['h0991]=8'h09; mem['h0992]=8'h3A; mem['h0993]=8'h2C;
    mem['h0994]=8'h81; mem['h0995]=8'hFE; mem['h0996]=8'h90; mem['h0997]=8'hDA;
    mem['h0998]=8'hD7; mem['h0999]=8'h17; mem['h099A]=8'h01; mem['h099B]=8'h80;
    mem['h099C]=8'h90; mem['h099D]=8'h11; mem['h099E]=8'h00; mem['h099F]=8'h00;
    mem['h09A0]=8'hE5; mem['h09A1]=8'hCD; mem['h09A2]=8'hAA; mem['h09A3]=8'h17;
    mem['h09A4]=8'hE1; mem['h09A5]=8'h51; mem['h09A6]=8'hC8; mem['h09A7]=8'h1E;
    mem['h09A8]=8'h08; mem['h09A9]=8'hC3; mem['h09AA]=8'h9C; mem['h09AB]=8'h04;
    mem['h09AC]=8'h2B; mem['h09AD]=8'h11; mem['h09AE]=8'h00; mem['h09AF]=8'h00;
    mem['h09B0]=8'hCD; mem['h09B1]=8'hE0; mem['h09B2]=8'h08; mem['h09B3]=8'hD0;
    mem['h09B4]=8'hE5; mem['h09B5]=8'hF5; mem['h09B6]=8'h21; mem['h09B7]=8'h98;
    mem['h09B8]=8'h19; mem['h09B9]=8'hCD; mem['h09BA]=8'h50; mem['h09BB]=8'h07;
    mem['h09BC]=8'hDA; mem['h09BD]=8'h88; mem['h09BE]=8'h04; mem['h09BF]=8'h62;
    mem['h09C0]=8'h6B; mem['h09C1]=8'h19; mem['h09C2]=8'h29; mem['h09C3]=8'h19;
    mem['h09C4]=8'h29; mem['h09C5]=8'hF1; mem['h09C6]=8'hD6; mem['h09C7]=8'h30;
    mem['h09C8]=8'h5F; mem['h09C9]=8'h16; mem['h09CA]=8'h00; mem['h09CB]=8'h19;
    mem['h09CC]=8'hEB; mem['h09CD]=8'hE1; mem['h09CE]=8'hC3; mem['h09CF]=8'hB0;
    mem['h09D0]=8'h09; mem['h09D1]=8'hCA; mem['h09D2]=8'hA4; mem['h09D3]=8'h05;
    mem['h09D4]=8'hCD; mem['h09D5]=8'h89; mem['h09D6]=8'h09; mem['h09D7]=8'h2B;
    mem['h09D8]=8'hCD; mem['h09D9]=8'hE0; mem['h09DA]=8'h08; mem['h09DB]=8'hE5;
    mem['h09DC]=8'h2A; mem['h09DD]=8'hF4; mem['h09DE]=8'h80; mem['h09DF]=8'hCA;
    mem['h09E0]=8'hF4; mem['h09E1]=8'h09; mem['h09E2]=8'hE1; mem['h09E3]=8'hCD;
    mem['h09E4]=8'h56; mem['h09E5]=8'h07; mem['h09E6]=8'h2C; mem['h09E7]=8'hD5;
    mem['h09E8]=8'hCD; mem['h09E9]=8'h89; mem['h09EA]=8'h09; mem['h09EB]=8'h2B;
    mem['h09EC]=8'hCD; mem['h09ED]=8'hE0; mem['h09EE]=8'h08; mem['h09EF]=8'hC2;
    mem['h09F0]=8'h88; mem['h09F1]=8'h04; mem['h09F2]=8'hE3; mem['h09F3]=8'hEB;
    mem['h09F4]=8'h7D; mem['h09F5]=8'h93; mem['h09F6]=8'h5F; mem['h09F7]=8'h7C;
    mem['h09F8]=8'h9A; mem['h09F9]=8'h57; mem['h09FA]=8'hDA; mem['h09FB]=8'h7D;
    mem['h09FC]=8'h04; mem['h09FD]=8'hE5; mem['h09FE]=8'h2A; mem['h09FF]=8'h1B;
    mem['h0A00]=8'h81; mem['h0A01]=8'h01; mem['h0A02]=8'h28; mem['h0A03]=8'h00;
    mem['h0A04]=8'h09; mem['h0A05]=8'hCD; mem['h0A06]=8'h50; mem['h0A07]=8'h07;
    mem['h0A08]=8'hD2; mem['h0A09]=8'h7D; mem['h0A0A]=8'h04; mem['h0A0B]=8'hEB;
    mem['h0A0C]=8'h22; mem['h0A0D]=8'h9F; mem['h0A0E]=8'h80; mem['h0A0F]=8'hE1;
    mem['h0A10]=8'h22; mem['h0A11]=8'hF4; mem['h0A12]=8'h80; mem['h0A13]=8'hE1;
    mem['h0A14]=8'hC3; mem['h0A15]=8'hA4; mem['h0A16]=8'h05; mem['h0A17]=8'hCA;
    mem['h0A18]=8'hA0; mem['h0A19]=8'h05; mem['h0A1A]=8'hCD; mem['h0A1B]=8'hA4;
    mem['h0A1C]=8'h05; mem['h0A1D]=8'h01; mem['h0A1E]=8'hA0; mem['h0A1F]=8'h08;
    mem['h0A20]=8'hC3; mem['h0A21]=8'h33; mem['h0A22]=8'h0A; mem['h0A23]=8'h0E;
    mem['h0A24]=8'h03; mem['h0A25]=8'hCD; mem['h0A26]=8'h65; mem['h0A27]=8'h04;
    mem['h0A28]=8'hC1; mem['h0A29]=8'hE5; mem['h0A2A]=8'hE5; mem['h0A2B]=8'h2A;
    mem['h0A2C]=8'hA1; mem['h0A2D]=8'h80; mem['h0A2E]=8'hE3; mem['h0A2F]=8'h3E;
    mem['h0A30]=8'h8C; mem['h0A31]=8'hF5; mem['h0A32]=8'h33; mem['h0A33]=8'hC5;
    mem['h0A34]=8'hCD; mem['h0A35]=8'hAC; mem['h0A36]=8'h09; mem['h0A37]=8'hCD;
    mem['h0A38]=8'h79; mem['h0A39]=8'h0A; mem['h0A3A]=8'hE5; mem['h0A3B]=8'h2A;
    mem['h0A3C]=8'hA1; mem['h0A3D]=8'h80; mem['h0A3E]=8'hCD; mem['h0A3F]=8'h50;
    mem['h0A40]=8'h07; mem['h0A41]=8'hE1; mem['h0A42]=8'h23; mem['h0A43]=8'hDC;
    mem['h0A44]=8'h77; mem['h0A45]=8'h05; mem['h0A46]=8'hD4; mem['h0A47]=8'h74;
    mem['h0A48]=8'h05; mem['h0A49]=8'h60; mem['h0A4A]=8'h69; mem['h0A4B]=8'h2B;
    mem['h0A4C]=8'hD8; mem['h0A4D]=8'h1E; mem['h0A4E]=8'h0E; mem['h0A4F]=8'hC3;
    mem['h0A50]=8'h9C; mem['h0A51]=8'h04; mem['h0A52]=8'hC0; mem['h0A53]=8'h16;
    mem['h0A54]=8'hFF; mem['h0A55]=8'hCD; mem['h0A56]=8'h31; mem['h0A57]=8'h04;
    mem['h0A58]=8'hF9; mem['h0A59]=8'hFE; mem['h0A5A]=8'h8C; mem['h0A5B]=8'h1E;
    mem['h0A5C]=8'h04; mem['h0A5D]=8'hC2; mem['h0A5E]=8'h9C; mem['h0A5F]=8'h04;
    mem['h0A60]=8'hE1; mem['h0A61]=8'h22; mem['h0A62]=8'hA1; mem['h0A63]=8'h80;
    mem['h0A64]=8'h23; mem['h0A65]=8'h7C; mem['h0A66]=8'hB5; mem['h0A67]=8'hC2;
    mem['h0A68]=8'h71; mem['h0A69]=8'h0A; mem['h0A6A]=8'h3A; mem['h0A6B]=8'h11;
    mem['h0A6C]=8'h81; mem['h0A6D]=8'hB7; mem['h0A6E]=8'hC2; mem['h0A6F]=8'hD2;
    mem['h0A70]=8'h04; mem['h0A71]=8'h21; mem['h0A72]=8'hA0; mem['h0A73]=8'h08;
    mem['h0A74]=8'hE3; mem['h0A75]=8'h3E; mem['h0A76]=8'hE1; mem['h0A77]=8'h01;
    mem['h0A78]=8'h3A; mem['h0A79]=8'h0E; mem['h0A7A]=8'h00; mem['h0A7B]=8'h06;
    mem['h0A7C]=8'h00; mem['h0A7D]=8'h79; mem['h0A7E]=8'h48; mem['h0A7F]=8'h47;
    mem['h0A80]=8'h7E; mem['h0A81]=8'hB7; mem['h0A82]=8'hC8; mem['h0A83]=8'hB8;
    mem['h0A84]=8'hC8; mem['h0A85]=8'h23; mem['h0A86]=8'hFE; mem['h0A87]=8'h22;
    mem['h0A88]=8'hCA; mem['h0A89]=8'h7D; mem['h0A8A]=8'h0A; mem['h0A8B]=8'hC3;
    mem['h0A8C]=8'h80; mem['h0A8D]=8'h0A; mem['h0A8E]=8'hCD; mem['h0A8F]=8'h43;
    mem['h0A90]=8'h0F; mem['h0A91]=8'hCD; mem['h0A92]=8'h56; mem['h0A93]=8'h07;
    mem['h0A94]=8'hB4; mem['h0A95]=8'hD5; mem['h0A96]=8'h3A; mem['h0A97]=8'hF2;
    mem['h0A98]=8'h80; mem['h0A99]=8'hF5; mem['h0A9A]=8'hCD; mem['h0A9B]=8'h5F;
    mem['h0A9C]=8'h0D; mem['h0A9D]=8'hF1; mem['h0A9E]=8'hE3; mem['h0A9F]=8'h22;
    mem['h0AA0]=8'h13; mem['h0AA1]=8'h81; mem['h0AA2]=8'h1F; mem['h0AA3]=8'hCD;
    mem['h0AA4]=8'h52; mem['h0AA5]=8'h0D; mem['h0AA6]=8'hCA; mem['h0AA7]=8'hE1;
    mem['h0AA8]=8'h0A; mem['h0AA9]=8'hE5; mem['h0AAA]=8'h2A; mem['h0AAB]=8'h29;
    mem['h0AAC]=8'h81; mem['h0AAD]=8'hE5; mem['h0AAE]=8'h23; mem['h0AAF]=8'h23;
    mem['h0AB0]=8'h5E; mem['h0AB1]=8'h23; mem['h0AB2]=8'h56; mem['h0AB3]=8'h2A;
    mem['h0AB4]=8'hA3; mem['h0AB5]=8'h80; mem['h0AB6]=8'hCD; mem['h0AB7]=8'h50;
    mem['h0AB8]=8'h07; mem['h0AB9]=8'hD2; mem['h0ABA]=8'hD0; mem['h0ABB]=8'h0A;
    mem['h0ABC]=8'h2A; mem['h0ABD]=8'h9F; mem['h0ABE]=8'h80; mem['h0ABF]=8'hCD;
    mem['h0AC0]=8'h50; mem['h0AC1]=8'h07; mem['h0AC2]=8'hD1; mem['h0AC3]=8'hD2;
    mem['h0AC4]=8'hD8; mem['h0AC5]=8'h0A; mem['h0AC6]=8'h21; mem['h0AC7]=8'h04;
    mem['h0AC8]=8'h81; mem['h0AC9]=8'hCD; mem['h0ACA]=8'h50; mem['h0ACB]=8'h07;
    mem['h0ACC]=8'hD2; mem['h0ACD]=8'hD8; mem['h0ACE]=8'h0A; mem['h0ACF]=8'h3E;
    mem['h0AD0]=8'hD1; mem['h0AD1]=8'hCD; mem['h0AD2]=8'h87; mem['h0AD3]=8'h13;
    mem['h0AD4]=8'hEB; mem['h0AD5]=8'hCD; mem['h0AD6]=8'hC0; mem['h0AD7]=8'h11;
    mem['h0AD8]=8'hCD; mem['h0AD9]=8'h87; mem['h0ADA]=8'h13; mem['h0ADB]=8'hE1;
    mem['h0ADC]=8'hCD; mem['h0ADD]=8'h8A; mem['h0ADE]=8'h17; mem['h0ADF]=8'hE1;
    mem['h0AE0]=8'hC9; mem['h0AE1]=8'hE5; mem['h0AE2]=8'hCD; mem['h0AE3]=8'h87;
    mem['h0AE4]=8'h17; mem['h0AE5]=8'hD1; mem['h0AE6]=8'hE1; mem['h0AE7]=8'hC9;
    mem['h0AE8]=8'hCD; mem['h0AE9]=8'hAE; mem['h0AEA]=8'h14; mem['h0AEB]=8'h7E;
    mem['h0AEC]=8'h47; mem['h0AED]=8'hFE; mem['h0AEE]=8'h8C; mem['h0AEF]=8'hCA;
    mem['h0AF0]=8'hF7; mem['h0AF1]=8'h0A; mem['h0AF2]=8'hCD; mem['h0AF3]=8'h56;
    mem['h0AF4]=8'h07; mem['h0AF5]=8'h88; mem['h0AF6]=8'h2B; mem['h0AF7]=8'h4B;
    mem['h0AF8]=8'h0D; mem['h0AF9]=8'h78; mem['h0AFA]=8'hCA; mem['h0AFB]=8'hC8;
    mem['h0AFC]=8'h08; mem['h0AFD]=8'hCD; mem['h0AFE]=8'hAD; mem['h0AFF]=8'h09;
    mem['h0B00]=8'hFE; mem['h0B01]=8'h2C; mem['h0B02]=8'hC0; mem['h0B03]=8'hC3;
    mem['h0B04]=8'hF8; mem['h0B05]=8'h0A; mem['h0B06]=8'hCD; mem['h0B07]=8'h5F;
    mem['h0B08]=8'h0D; mem['h0B09]=8'h7E; mem['h0B0A]=8'hFE; mem['h0B0B]=8'h88;
    mem['h0B0C]=8'hCA; mem['h0B0D]=8'h14; mem['h0B0E]=8'h0B; mem['h0B0F]=8'hCD;
    mem['h0B10]=8'h56; mem['h0B11]=8'h07; mem['h0B12]=8'hA9; mem['h0B13]=8'h2B;
    mem['h0B14]=8'hCD; mem['h0B15]=8'h50; mem['h0B16]=8'h0D; mem['h0B17]=8'hCD;
    mem['h0B18]=8'h2F; mem['h0B19]=8'h17; mem['h0B1A]=8'hCA; mem['h0B1B]=8'h79;
    mem['h0B1C]=8'h0A; mem['h0B1D]=8'hCD; mem['h0B1E]=8'hE0; mem['h0B1F]=8'h08;
    mem['h0B20]=8'hDA; mem['h0B21]=8'h34; mem['h0B22]=8'h0A; mem['h0B23]=8'hC3;
    mem['h0B24]=8'hC7; mem['h0B25]=8'h08; mem['h0B26]=8'h2B; mem['h0B27]=8'hCD;
    mem['h0B28]=8'hE0; mem['h0B29]=8'h08; mem['h0B2A]=8'hCA; mem['h0B2B]=8'h88;
    mem['h0B2C]=8'h0B; mem['h0B2D]=8'hC8; mem['h0B2E]=8'hFE; mem['h0B2F]=8'hA5;
    mem['h0B30]=8'hCA; mem['h0B31]=8'hBB; mem['h0B32]=8'h0B; mem['h0B33]=8'hFE;
    mem['h0B34]=8'hA8; mem['h0B35]=8'hCA; mem['h0B36]=8'hBB; mem['h0B37]=8'h0B;
    mem['h0B38]=8'hE5; mem['h0B39]=8'hFE; mem['h0B3A]=8'h2C; mem['h0B3B]=8'hCA;
    mem['h0B3C]=8'hA4; mem['h0B3D]=8'h0B; mem['h0B3E]=8'hFE; mem['h0B3F]=8'h3B;
    mem['h0B40]=8'hCA; mem['h0B41]=8'hDE; mem['h0B42]=8'h0B; mem['h0B43]=8'hC1;
    mem['h0B44]=8'hCD; mem['h0B45]=8'h5F; mem['h0B46]=8'h0D; mem['h0B47]=8'hE5;
    mem['h0B48]=8'h3A; mem['h0B49]=8'hF2; mem['h0B4A]=8'h80; mem['h0B4B]=8'hB7;
    mem['h0B4C]=8'hC2; mem['h0B4D]=8'h74; mem['h0B4E]=8'h0B; mem['h0B4F]=8'hCD;
    mem['h0B50]=8'hD4; mem['h0B51]=8'h18; mem['h0B52]=8'hCD; mem['h0B53]=8'hE4;
    mem['h0B54]=8'h11; mem['h0B55]=8'h36; mem['h0B56]=8'h20; mem['h0B57]=8'h2A;
    mem['h0B58]=8'h29; mem['h0B59]=8'h81; mem['h0B5A]=8'h34; mem['h0B5B]=8'h2A;
    mem['h0B5C]=8'h29; mem['h0B5D]=8'h81; mem['h0B5E]=8'h3A; mem['h0B5F]=8'h87;
    mem['h0B60]=8'h80; mem['h0B61]=8'h47; mem['h0B62]=8'h04; mem['h0B63]=8'hCA;
    mem['h0B64]=8'h70; mem['h0B65]=8'h0B; mem['h0B66]=8'h04; mem['h0B67]=8'h3A;
    mem['h0B68]=8'hF0; mem['h0B69]=8'h80; mem['h0B6A]=8'h86; mem['h0B6B]=8'h3D;
    mem['h0B6C]=8'hB8; mem['h0B6D]=8'hD4; mem['h0B6E]=8'h88; mem['h0B6F]=8'h0B;
    mem['h0B70]=8'hCD; mem['h0B71]=8'h29; mem['h0B72]=8'h12; mem['h0B73]=8'hAF;
    mem['h0B74]=8'hC4; mem['h0B75]=8'h29; mem['h0B76]=8'h12; mem['h0B77]=8'hE1;
    mem['h0B78]=8'hC3; mem['h0B79]=8'h26; mem['h0B7A]=8'h0B; mem['h0B7B]=8'h3A;
    mem['h0B7C]=8'hF0; mem['h0B7D]=8'h80; mem['h0B7E]=8'hB7; mem['h0B7F]=8'hC8;
    mem['h0B80]=8'hC3; mem['h0B81]=8'h88; mem['h0B82]=8'h0B; mem['h0B83]=8'h36;
    mem['h0B84]=8'h00; mem['h0B85]=8'h21; mem['h0B86]=8'hA5; mem['h0B87]=8'h80;
    mem['h0B88]=8'h3E; mem['h0B89]=8'h0D; mem['h0B8A]=8'hCD; mem['h0B8B]=8'h61;
    mem['h0B8C]=8'h07; mem['h0B8D]=8'h3E; mem['h0B8E]=8'h0A; mem['h0B8F]=8'hCD;
    mem['h0B90]=8'h61; mem['h0B91]=8'h07; mem['h0B92]=8'hAF; mem['h0B93]=8'h32;
    mem['h0B94]=8'hF0; mem['h0B95]=8'h80; mem['h0B96]=8'h3A; mem['h0B97]=8'h86;
    mem['h0B98]=8'h80; mem['h0B99]=8'h3D; mem['h0B9A]=8'hC8; mem['h0B9B]=8'hF5;
    mem['h0B9C]=8'hAF; mem['h0B9D]=8'hCD; mem['h0B9E]=8'h61; mem['h0B9F]=8'h07;
    mem['h0BA0]=8'hF1; mem['h0BA1]=8'hC3; mem['h0BA2]=8'h99; mem['h0BA3]=8'h0B;
    mem['h0BA4]=8'h3A; mem['h0BA5]=8'h88; mem['h0BA6]=8'h80; mem['h0BA7]=8'h47;
    mem['h0BA8]=8'h3A; mem['h0BA9]=8'hF0; mem['h0BAA]=8'h80; mem['h0BAB]=8'hB8;
    mem['h0BAC]=8'hD4; mem['h0BAD]=8'h88; mem['h0BAE]=8'h0B; mem['h0BAF]=8'hD2;
    mem['h0BB0]=8'hDE; mem['h0BB1]=8'h0B; mem['h0BB2]=8'hD6; mem['h0BB3]=8'h0E;
    mem['h0BB4]=8'hD2; mem['h0BB5]=8'hB2; mem['h0BB6]=8'h0B; mem['h0BB7]=8'h2F;
    mem['h0BB8]=8'hC3; mem['h0BB9]=8'hD3; mem['h0BBA]=8'h0B; mem['h0BBB]=8'hF5;
    mem['h0BBC]=8'hCD; mem['h0BBD]=8'hAB; mem['h0BBE]=8'h14; mem['h0BBF]=8'hCD;
    mem['h0BC0]=8'h56; mem['h0BC1]=8'h07; mem['h0BC2]=8'h29; mem['h0BC3]=8'h2B;
    mem['h0BC4]=8'hF1; mem['h0BC5]=8'hD6; mem['h0BC6]=8'hA8; mem['h0BC7]=8'hE5;
    mem['h0BC8]=8'hCA; mem['h0BC9]=8'hCE; mem['h0BCA]=8'h0B; mem['h0BCB]=8'h3A;
    mem['h0BCC]=8'hF0; mem['h0BCD]=8'h80; mem['h0BCE]=8'h2F; mem['h0BCF]=8'h83;
    mem['h0BD0]=8'hD2; mem['h0BD1]=8'hDE; mem['h0BD2]=8'h0B; mem['h0BD3]=8'h3C;
    mem['h0BD4]=8'h47; mem['h0BD5]=8'h3E; mem['h0BD6]=8'h20; mem['h0BD7]=8'hCD;
    mem['h0BD8]=8'h61; mem['h0BD9]=8'h07; mem['h0BDA]=8'h05; mem['h0BDB]=8'hC2;
    mem['h0BDC]=8'hD7; mem['h0BDD]=8'h0B; mem['h0BDE]=8'hE1; mem['h0BDF]=8'hCD;
    mem['h0BE0]=8'hE0; mem['h0BE1]=8'h08; mem['h0BE2]=8'hC3; mem['h0BE3]=8'h2D;
    mem['h0BE4]=8'h0B; mem['h0BE5]=8'h3F; mem['h0BE6]=8'h52; mem['h0BE7]=8'h65;
    mem['h0BE8]=8'h64; mem['h0BE9]=8'h6F; mem['h0BEA]=8'h20; mem['h0BEB]=8'h66;
    mem['h0BEC]=8'h72; mem['h0BED]=8'h6F; mem['h0BEE]=8'h6D; mem['h0BEF]=8'h20;
    mem['h0BF0]=8'h73; mem['h0BF1]=8'h74; mem['h0BF2]=8'h61; mem['h0BF3]=8'h72;
    mem['h0BF4]=8'h74; mem['h0BF5]=8'h0D; mem['h0BF6]=8'h0A; mem['h0BF7]=8'h00;
    mem['h0BF8]=8'h3A; mem['h0BF9]=8'h12; mem['h0BFA]=8'h81; mem['h0BFB]=8'hB7;
    mem['h0BFC]=8'hC2; mem['h0BFD]=8'h82; mem['h0BFE]=8'h04; mem['h0BFF]=8'hC1;
    mem['h0C00]=8'h21; mem['h0C01]=8'hE5; mem['h0C02]=8'h0B; mem['h0C03]=8'hCD;
    mem['h0C04]=8'h26; mem['h0C05]=8'h12; mem['h0C06]=8'hC3; mem['h0C07]=8'hD3;
    mem['h0C08]=8'h05; mem['h0C09]=8'hCD; mem['h0C0A]=8'h91; mem['h0C0B]=8'h11;
    mem['h0C0C]=8'h7E; mem['h0C0D]=8'hFE; mem['h0C0E]=8'h22; mem['h0C0F]=8'h3E;
    mem['h0C10]=8'h00; mem['h0C11]=8'h32; mem['h0C12]=8'h8A; mem['h0C13]=8'h80;
    mem['h0C14]=8'hC2; mem['h0C15]=8'h23; mem['h0C16]=8'h0C; mem['h0C17]=8'hCD;
    mem['h0C18]=8'hE5; mem['h0C19]=8'h11; mem['h0C1A]=8'hCD; mem['h0C1B]=8'h56;
    mem['h0C1C]=8'h07; mem['h0C1D]=8'h3B; mem['h0C1E]=8'hE5; mem['h0C1F]=8'hCD;
    mem['h0C20]=8'h29; mem['h0C21]=8'h12; mem['h0C22]=8'h3E; mem['h0C23]=8'hE5;
    mem['h0C24]=8'hCD; mem['h0C25]=8'hD7; mem['h0C26]=8'h05; mem['h0C27]=8'hC1;
    mem['h0C28]=8'hDA; mem['h0C29]=8'h2F; mem['h0C2A]=8'h09; mem['h0C2B]=8'h23;
    mem['h0C2C]=8'h7E; mem['h0C2D]=8'hB7; mem['h0C2E]=8'h2B; mem['h0C2F]=8'hC5;
    mem['h0C30]=8'hCA; mem['h0C31]=8'h76; mem['h0C32]=8'h0A; mem['h0C33]=8'h36;
    mem['h0C34]=8'h2C; mem['h0C35]=8'hC3; mem['h0C36]=8'h3D; mem['h0C37]=8'h0C;
    mem['h0C38]=8'hE5; mem['h0C39]=8'h2A; mem['h0C3A]=8'h21; mem['h0C3B]=8'h81;
    mem['h0C3C]=8'hF6; mem['h0C3D]=8'hAF; mem['h0C3E]=8'h32; mem['h0C3F]=8'h12;
    mem['h0C40]=8'h81; mem['h0C41]=8'hE3; mem['h0C42]=8'hC3; mem['h0C43]=8'h49;
    mem['h0C44]=8'h0C; mem['h0C45]=8'hCD; mem['h0C46]=8'h56; mem['h0C47]=8'h07;
    mem['h0C48]=8'h2C; mem['h0C49]=8'hCD; mem['h0C4A]=8'h43; mem['h0C4B]=8'h0F;
    mem['h0C4C]=8'hE3; mem['h0C4D]=8'hD5; mem['h0C4E]=8'h7E; mem['h0C4F]=8'hFE;
    mem['h0C50]=8'h2C; mem['h0C51]=8'hCA; mem['h0C52]=8'h71; mem['h0C53]=8'h0C;
    mem['h0C54]=8'h3A; mem['h0C55]=8'h12; mem['h0C56]=8'h81; mem['h0C57]=8'hB7;
    mem['h0C58]=8'hC2; mem['h0C59]=8'hDE; mem['h0C5A]=8'h0C; mem['h0C5B]=8'h3E;
    mem['h0C5C]=8'h3F; mem['h0C5D]=8'hCD; mem['h0C5E]=8'h61; mem['h0C5F]=8'h07;
    mem['h0C60]=8'hCD; mem['h0C61]=8'hD7; mem['h0C62]=8'h05; mem['h0C63]=8'hD1;
    mem['h0C64]=8'hC1; mem['h0C65]=8'hDA; mem['h0C66]=8'h2F; mem['h0C67]=8'h09;
    mem['h0C68]=8'h23; mem['h0C69]=8'h7E; mem['h0C6A]=8'hB7; mem['h0C6B]=8'h2B;
    mem['h0C6C]=8'hC5; mem['h0C6D]=8'hCA; mem['h0C6E]=8'h76; mem['h0C6F]=8'h0A;
    mem['h0C70]=8'hD5; mem['h0C71]=8'h3A; mem['h0C72]=8'hF2; mem['h0C73]=8'h80;
    mem['h0C74]=8'hB7; mem['h0C75]=8'hCA; mem['h0C76]=8'h9B; mem['h0C77]=8'h0C;
    mem['h0C78]=8'hCD; mem['h0C79]=8'hE0; mem['h0C7A]=8'h08; mem['h0C7B]=8'h57;
    mem['h0C7C]=8'h47; mem['h0C7D]=8'hFE; mem['h0C7E]=8'h22; mem['h0C7F]=8'hCA;
    mem['h0C80]=8'h8F; mem['h0C81]=8'h0C; mem['h0C82]=8'h3A; mem['h0C83]=8'h12;
    mem['h0C84]=8'h81; mem['h0C85]=8'hB7; mem['h0C86]=8'h57; mem['h0C87]=8'hCA;
    mem['h0C88]=8'h8C; mem['h0C89]=8'h0C; mem['h0C8A]=8'h16; mem['h0C8B]=8'h3A;
    mem['h0C8C]=8'h06; mem['h0C8D]=8'h2C; mem['h0C8E]=8'h2B; mem['h0C8F]=8'hCD;
    mem['h0C90]=8'hE8; mem['h0C91]=8'h11; mem['h0C92]=8'hEB; mem['h0C93]=8'h21;
    mem['h0C94]=8'hA6; mem['h0C95]=8'h0C; mem['h0C96]=8'hE3; mem['h0C97]=8'hD5;
    mem['h0C98]=8'hC3; mem['h0C99]=8'hA9; mem['h0C9A]=8'h0A; mem['h0C9B]=8'hCD;
    mem['h0C9C]=8'hE0; mem['h0C9D]=8'h08; mem['h0C9E]=8'hCD; mem['h0C9F]=8'h36;
    mem['h0CA0]=8'h18; mem['h0CA1]=8'hE3; mem['h0CA2]=8'hCD; mem['h0CA3]=8'h87;
    mem['h0CA4]=8'h17; mem['h0CA5]=8'hE1; mem['h0CA6]=8'h2B; mem['h0CA7]=8'hCD;
    mem['h0CA8]=8'hE0; mem['h0CA9]=8'h08; mem['h0CAA]=8'hCA; mem['h0CAB]=8'hB2;
    mem['h0CAC]=8'h0C; mem['h0CAD]=8'hFE; mem['h0CAE]=8'h2C; mem['h0CAF]=8'hC2;
    mem['h0CB0]=8'hF8; mem['h0CB1]=8'h0B; mem['h0CB2]=8'hE3; mem['h0CB3]=8'h2B;
    mem['h0CB4]=8'hCD; mem['h0CB5]=8'hE0; mem['h0CB6]=8'h08; mem['h0CB7]=8'hC2;
    mem['h0CB8]=8'h45; mem['h0CB9]=8'h0C; mem['h0CBA]=8'hD1; mem['h0CBB]=8'h3A;
    mem['h0CBC]=8'h12; mem['h0CBD]=8'h81; mem['h0CBE]=8'hB7; mem['h0CBF]=8'hEB;
    mem['h0CC0]=8'hC2; mem['h0CC1]=8'h06; mem['h0CC2]=8'h09; mem['h0CC3]=8'hD5;
    mem['h0CC4]=8'hB6; mem['h0CC5]=8'h21; mem['h0CC6]=8'hCD; mem['h0CC7]=8'h0C;
    mem['h0CC8]=8'hC4; mem['h0CC9]=8'h26; mem['h0CCA]=8'h12; mem['h0CCB]=8'hE1;
    mem['h0CCC]=8'hC9; mem['h0CCD]=8'h3F; mem['h0CCE]=8'h45; mem['h0CCF]=8'h78;
    mem['h0CD0]=8'h74; mem['h0CD1]=8'h72; mem['h0CD2]=8'h61; mem['h0CD3]=8'h20;
    mem['h0CD4]=8'h69; mem['h0CD5]=8'h67; mem['h0CD6]=8'h6E; mem['h0CD7]=8'h6F;
    mem['h0CD8]=8'h72; mem['h0CD9]=8'h65; mem['h0CDA]=8'h64; mem['h0CDB]=8'h0D;
    mem['h0CDC]=8'h0A; mem['h0CDD]=8'h00; mem['h0CDE]=8'hCD; mem['h0CDF]=8'h77;
    mem['h0CE0]=8'h0A; mem['h0CE1]=8'hB7; mem['h0CE2]=8'hC2; mem['h0CE3]=8'hF7;
    mem['h0CE4]=8'h0C; mem['h0CE5]=8'h23; mem['h0CE6]=8'h7E; mem['h0CE7]=8'h23;
    mem['h0CE8]=8'hB6; mem['h0CE9]=8'h1E; mem['h0CEA]=8'h06; mem['h0CEB]=8'hCA;
    mem['h0CEC]=8'h9C; mem['h0CED]=8'h04; mem['h0CEE]=8'h23; mem['h0CEF]=8'h5E;
    mem['h0CF0]=8'h23; mem['h0CF1]=8'h56; mem['h0CF2]=8'hEB; mem['h0CF3]=8'h22;
    mem['h0CF4]=8'h0E; mem['h0CF5]=8'h81; mem['h0CF6]=8'hEB; mem['h0CF7]=8'hCD;
    mem['h0CF8]=8'hE0; mem['h0CF9]=8'h08; mem['h0CFA]=8'hFE; mem['h0CFB]=8'h83;
    mem['h0CFC]=8'hC2; mem['h0CFD]=8'hDE; mem['h0CFE]=8'h0C; mem['h0CFF]=8'hC3;
    mem['h0D00]=8'h71; mem['h0D01]=8'h0C; mem['h0D02]=8'h11; mem['h0D03]=8'h00;
    mem['h0D04]=8'h00; mem['h0D05]=8'hC4; mem['h0D06]=8'h43; mem['h0D07]=8'h0F;
    mem['h0D08]=8'h22; mem['h0D09]=8'h13; mem['h0D0A]=8'h81; mem['h0D0B]=8'hCD;
    mem['h0D0C]=8'h31; mem['h0D0D]=8'h04; mem['h0D0E]=8'hC2; mem['h0D0F]=8'h8E;
    mem['h0D10]=8'h04; mem['h0D11]=8'hF9; mem['h0D12]=8'hD5; mem['h0D13]=8'h7E;
    mem['h0D14]=8'h23; mem['h0D15]=8'hF5; mem['h0D16]=8'hD5; mem['h0D17]=8'hCD;
    mem['h0D18]=8'h6D; mem['h0D19]=8'h17; mem['h0D1A]=8'hE3; mem['h0D1B]=8'hE5;
    mem['h0D1C]=8'hCD; mem['h0D1D]=8'hDA; mem['h0D1E]=8'h14; mem['h0D1F]=8'hE1;
    mem['h0D20]=8'hCD; mem['h0D21]=8'h87; mem['h0D22]=8'h17; mem['h0D23]=8'hE1;
    mem['h0D24]=8'hCD; mem['h0D25]=8'h7E; mem['h0D26]=8'h17; mem['h0D27]=8'hE5;
    mem['h0D28]=8'hCD; mem['h0D29]=8'hAA; mem['h0D2A]=8'h17; mem['h0D2B]=8'hE1;
    mem['h0D2C]=8'hC1; mem['h0D2D]=8'h90; mem['h0D2E]=8'hCD; mem['h0D2F]=8'h7E;
    mem['h0D30]=8'h17; mem['h0D31]=8'hCA; mem['h0D32]=8'h3D; mem['h0D33]=8'h0D;
    mem['h0D34]=8'hEB; mem['h0D35]=8'h22; mem['h0D36]=8'hA1; mem['h0D37]=8'h80;
    mem['h0D38]=8'h69; mem['h0D39]=8'h60; mem['h0D3A]=8'hC3; mem['h0D3B]=8'h9C;
    mem['h0D3C]=8'h08; mem['h0D3D]=8'hF9; mem['h0D3E]=8'h2A; mem['h0D3F]=8'h13;
    mem['h0D40]=8'h81; mem['h0D41]=8'h7E; mem['h0D42]=8'hFE; mem['h0D43]=8'h2C;
    mem['h0D44]=8'hC2; mem['h0D45]=8'hA0; mem['h0D46]=8'h08; mem['h0D47]=8'hCD;
    mem['h0D48]=8'hE0; mem['h0D49]=8'h08; mem['h0D4A]=8'hCD; mem['h0D4B]=8'h05;
    mem['h0D4C]=8'h0D; mem['h0D4D]=8'hCD; mem['h0D4E]=8'h5F; mem['h0D4F]=8'h0D;
    mem['h0D50]=8'hF6; mem['h0D51]=8'h37; mem['h0D52]=8'h3A; mem['h0D53]=8'hF2;
    mem['h0D54]=8'h80; mem['h0D55]=8'h8F; mem['h0D56]=8'hB7; mem['h0D57]=8'hE8;
    mem['h0D58]=8'hC3; mem['h0D59]=8'h9A; mem['h0D5A]=8'h04; mem['h0D5B]=8'hCD;
    mem['h0D5C]=8'h56; mem['h0D5D]=8'h07; mem['h0D5E]=8'h28; mem['h0D5F]=8'h2B;
    mem['h0D60]=8'h16; mem['h0D61]=8'h00; mem['h0D62]=8'hD5; mem['h0D63]=8'h0E;
    mem['h0D64]=8'h01; mem['h0D65]=8'hCD; mem['h0D66]=8'h65; mem['h0D67]=8'h04;
    mem['h0D68]=8'hCD; mem['h0D69]=8'hD6; mem['h0D6A]=8'h0D; mem['h0D6B]=8'h22;
    mem['h0D6C]=8'h15; mem['h0D6D]=8'h81; mem['h0D6E]=8'h2A; mem['h0D6F]=8'h15;
    mem['h0D70]=8'h81; mem['h0D71]=8'hC1; mem['h0D72]=8'h78; mem['h0D73]=8'hFE;
    mem['h0D74]=8'h78; mem['h0D75]=8'hD4; mem['h0D76]=8'h50; mem['h0D77]=8'h0D;
    mem['h0D78]=8'h7E; mem['h0D79]=8'h16; mem['h0D7A]=8'h00; mem['h0D7B]=8'hD6;
    mem['h0D7C]=8'hB3; mem['h0D7D]=8'hDA; mem['h0D7E]=8'h97; mem['h0D7F]=8'h0D;
    mem['h0D80]=8'hFE; mem['h0D81]=8'h03; mem['h0D82]=8'hD2; mem['h0D83]=8'h97;
    mem['h0D84]=8'h0D; mem['h0D85]=8'hFE; mem['h0D86]=8'h01; mem['h0D87]=8'h17;
    mem['h0D88]=8'hAA; mem['h0D89]=8'hBA; mem['h0D8A]=8'h57; mem['h0D8B]=8'hDA;
    mem['h0D8C]=8'h88; mem['h0D8D]=8'h04; mem['h0D8E]=8'h22; mem['h0D8F]=8'h0A;
    mem['h0D90]=8'h81; mem['h0D91]=8'hCD; mem['h0D92]=8'hE0; mem['h0D93]=8'h08;
    mem['h0D94]=8'hC3; mem['h0D95]=8'h7B; mem['h0D96]=8'h0D; mem['h0D97]=8'h7A;
    mem['h0D98]=8'hB7; mem['h0D99]=8'hC2; mem['h0D9A]=8'hBE; mem['h0D9B]=8'h0E;
    mem['h0D9C]=8'h7E; mem['h0D9D]=8'h22; mem['h0D9E]=8'h0A; mem['h0D9F]=8'h81;
    mem['h0DA0]=8'hD6; mem['h0DA1]=8'hAC; mem['h0DA2]=8'hD8; mem['h0DA3]=8'hFE;
    mem['h0DA4]=8'h07; mem['h0DA5]=8'hD0; mem['h0DA6]=8'h5F; mem['h0DA7]=8'h3A;
    mem['h0DA8]=8'hF2; mem['h0DA9]=8'h80; mem['h0DAA]=8'h3D; mem['h0DAB]=8'hB3;
    mem['h0DAC]=8'h7B; mem['h0DAD]=8'hCA; mem['h0DAE]=8'h1C; mem['h0DAF]=8'h13;
    mem['h0DB0]=8'h07; mem['h0DB1]=8'h83; mem['h0DB2]=8'h5F; mem['h0DB3]=8'h21;
    mem['h0DB4]=8'h7A; mem['h0DB5]=8'h03; mem['h0DB6]=8'h19; mem['h0DB7]=8'h78;
    mem['h0DB8]=8'h56; mem['h0DB9]=8'hBA; mem['h0DBA]=8'hD0; mem['h0DBB]=8'h23;
    mem['h0DBC]=8'hCD; mem['h0DBD]=8'h50; mem['h0DBE]=8'h0D; mem['h0DBF]=8'hC5;
    mem['h0DC0]=8'h01; mem['h0DC1]=8'h6E; mem['h0DC2]=8'h0D; mem['h0DC3]=8'hC5;
    mem['h0DC4]=8'h43; mem['h0DC5]=8'h4A; mem['h0DC6]=8'hCD; mem['h0DC7]=8'h60;
    mem['h0DC8]=8'h17; mem['h0DC9]=8'h58; mem['h0DCA]=8'h51; mem['h0DCB]=8'h4E;
    mem['h0DCC]=8'h23; mem['h0DCD]=8'h46; mem['h0DCE]=8'h23; mem['h0DCF]=8'hC5;
    mem['h0DD0]=8'h2A; mem['h0DD1]=8'h0A; mem['h0DD2]=8'h81; mem['h0DD3]=8'hC3;
    mem['h0DD4]=8'h62; mem['h0DD5]=8'h0D; mem['h0DD6]=8'hAF; mem['h0DD7]=8'h32;
    mem['h0DD8]=8'hF2; mem['h0DD9]=8'h80; mem['h0DDA]=8'hCD; mem['h0DDB]=8'hE0;
    mem['h0DDC]=8'h08; mem['h0DDD]=8'h1E; mem['h0DDE]=8'h24; mem['h0DDF]=8'hCA;
    mem['h0DE0]=8'h9C; mem['h0DE1]=8'h04; mem['h0DE2]=8'hDA; mem['h0DE3]=8'h36;
    mem['h0DE4]=8'h18; mem['h0DE5]=8'hCD; mem['h0DE6]=8'h7E; mem['h0DE7]=8'h09;
    mem['h0DE8]=8'hD2; mem['h0DE9]=8'h3D; mem['h0DEA]=8'h0E; mem['h0DEB]=8'hFE;
    mem['h0DEC]=8'h26; mem['h0DED]=8'h20; mem['h0DEE]=8'h12; mem['h0DEF]=8'hCD;
    mem['h0DF0]=8'hE0; mem['h0DF1]=8'h08; mem['h0DF2]=8'hFE; mem['h0DF3]=8'h48;
    mem['h0DF4]=8'hCA; mem['h0DF5]=8'h7A; mem['h0DF6]=8'h1C; mem['h0DF7]=8'hFE;
    mem['h0DF8]=8'h42; mem['h0DF9]=8'hCA; mem['h0DFA]=8'hEA; mem['h0DFB]=8'h1C;
    mem['h0DFC]=8'h1E; mem['h0DFD]=8'h02; mem['h0DFE]=8'hCA; mem['h0DFF]=8'h9C;
    mem['h0E00]=8'h04; mem['h0E01]=8'hFE; mem['h0E02]=8'hAC; mem['h0E03]=8'hCA;
    mem['h0E04]=8'hD6; mem['h0E05]=8'h0D; mem['h0E06]=8'hFE; mem['h0E07]=8'h2E;
    mem['h0E08]=8'hCA; mem['h0E09]=8'h36; mem['h0E0A]=8'h18; mem['h0E0B]=8'hFE;
    mem['h0E0C]=8'hAD; mem['h0E0D]=8'hCA; mem['h0E0E]=8'h2C; mem['h0E0F]=8'h0E;
    mem['h0E10]=8'hFE; mem['h0E11]=8'h22; mem['h0E12]=8'hCA; mem['h0E13]=8'hE5;
    mem['h0E14]=8'h11; mem['h0E15]=8'hFE; mem['h0E16]=8'hAA; mem['h0E17]=8'hCA;
    mem['h0E18]=8'h1E; mem['h0E19]=8'h0F; mem['h0E1A]=8'hFE; mem['h0E1B]=8'hA7;
    mem['h0E1C]=8'hCA; mem['h0E1D]=8'h49; mem['h0E1E]=8'h11; mem['h0E1F]=8'hD6;
    mem['h0E20]=8'hB6; mem['h0E21]=8'hD2; mem['h0E22]=8'h4E; mem['h0E23]=8'h0E;
    mem['h0E24]=8'hCD; mem['h0E25]=8'h5B; mem['h0E26]=8'h0D; mem['h0E27]=8'hCD;
    mem['h0E28]=8'h56; mem['h0E29]=8'h07; mem['h0E2A]=8'h29; mem['h0E2B]=8'hC9;
    mem['h0E2C]=8'h16; mem['h0E2D]=8'h7D; mem['h0E2E]=8'hCD; mem['h0E2F]=8'h62;
    mem['h0E30]=8'h0D; mem['h0E31]=8'h2A; mem['h0E32]=8'h15; mem['h0E33]=8'h81;
    mem['h0E34]=8'hE5; mem['h0E35]=8'hCD; mem['h0E36]=8'h58; mem['h0E37]=8'h17;
    mem['h0E38]=8'hCD; mem['h0E39]=8'h50; mem['h0E3A]=8'h0D; mem['h0E3B]=8'hE1;
    mem['h0E3C]=8'hC9; mem['h0E3D]=8'hCD; mem['h0E3E]=8'h43; mem['h0E3F]=8'h0F;
    mem['h0E40]=8'hE5; mem['h0E41]=8'hEB; mem['h0E42]=8'h22; mem['h0E43]=8'h29;
    mem['h0E44]=8'h81; mem['h0E45]=8'h3A; mem['h0E46]=8'hF2; mem['h0E47]=8'h80;
    mem['h0E48]=8'hB7; mem['h0E49]=8'hCC; mem['h0E4A]=8'h6D; mem['h0E4B]=8'h17;
    mem['h0E4C]=8'hE1; mem['h0E4D]=8'hC9; mem['h0E4E]=8'h06; mem['h0E4F]=8'h00;
    mem['h0E50]=8'h07; mem['h0E51]=8'h4F; mem['h0E52]=8'hC5; mem['h0E53]=8'hCD;
    mem['h0E54]=8'hE0; mem['h0E55]=8'h08; mem['h0E56]=8'h79; mem['h0E57]=8'hFE;
    mem['h0E58]=8'h31; mem['h0E59]=8'hDA; mem['h0E5A]=8'h75; mem['h0E5B]=8'h0E;
    mem['h0E5C]=8'hCD; mem['h0E5D]=8'h5B; mem['h0E5E]=8'h0D; mem['h0E5F]=8'hCD;
    mem['h0E60]=8'h56; mem['h0E61]=8'h07; mem['h0E62]=8'h2C; mem['h0E63]=8'hCD;
    mem['h0E64]=8'h51; mem['h0E65]=8'h0D; mem['h0E66]=8'hEB; mem['h0E67]=8'h2A;
    mem['h0E68]=8'h29; mem['h0E69]=8'h81; mem['h0E6A]=8'hE3; mem['h0E6B]=8'hE5;
    mem['h0E6C]=8'hEB; mem['h0E6D]=8'hCD; mem['h0E6E]=8'hAE; mem['h0E6F]=8'h14;
    mem['h0E70]=8'hEB; mem['h0E71]=8'hE3; mem['h0E72]=8'hC3; mem['h0E73]=8'h7D;
    mem['h0E74]=8'h0E; mem['h0E75]=8'hCD; mem['h0E76]=8'h24; mem['h0E77]=8'h0E;
    mem['h0E78]=8'hE3; mem['h0E79]=8'h11; mem['h0E7A]=8'h38; mem['h0E7B]=8'h0E;
    mem['h0E7C]=8'hD5; mem['h0E7D]=8'h01; mem['h0E7E]=8'hD9; mem['h0E7F]=8'h01;
    mem['h0E80]=8'h09; mem['h0E81]=8'h4E; mem['h0E82]=8'h23; mem['h0E83]=8'h66;
    mem['h0E84]=8'h69; mem['h0E85]=8'hE9; mem['h0E86]=8'h15; mem['h0E87]=8'hFE;
    mem['h0E88]=8'hAD; mem['h0E89]=8'hC8; mem['h0E8A]=8'hFE; mem['h0E8B]=8'h2D;
    mem['h0E8C]=8'hC8; mem['h0E8D]=8'h14; mem['h0E8E]=8'hFE; mem['h0E8F]=8'h2B;
    mem['h0E90]=8'hC8; mem['h0E91]=8'hFE; mem['h0E92]=8'hAC; mem['h0E93]=8'hC8;
    mem['h0E94]=8'h2B; mem['h0E95]=8'hC9; mem['h0E96]=8'hF6; mem['h0E97]=8'hAF;
    mem['h0E98]=8'hF5; mem['h0E99]=8'hCD; mem['h0E9A]=8'h50; mem['h0E9B]=8'h0D;
    mem['h0E9C]=8'hCD; mem['h0E9D]=8'h92; mem['h0E9E]=8'h09; mem['h0E9F]=8'hF1;
    mem['h0EA0]=8'hEB; mem['h0EA1]=8'hC1; mem['h0EA2]=8'hE3; mem['h0EA3]=8'hEB;
    mem['h0EA4]=8'hCD; mem['h0EA5]=8'h70; mem['h0EA6]=8'h17; mem['h0EA7]=8'hF5;
    mem['h0EA8]=8'hCD; mem['h0EA9]=8'h92; mem['h0EAA]=8'h09; mem['h0EAB]=8'hF1;
    mem['h0EAC]=8'hC1; mem['h0EAD]=8'h79; mem['h0EAE]=8'h21; mem['h0EAF]=8'h07;
    mem['h0EB0]=8'h11; mem['h0EB1]=8'hC2; mem['h0EB2]=8'hB9; mem['h0EB3]=8'h0E;
    mem['h0EB4]=8'hA3; mem['h0EB5]=8'h4F; mem['h0EB6]=8'h78; mem['h0EB7]=8'hA2;
    mem['h0EB8]=8'hE9; mem['h0EB9]=8'hB3; mem['h0EBA]=8'h4F; mem['h0EBB]=8'h78;
    mem['h0EBC]=8'hB2; mem['h0EBD]=8'hE9; mem['h0EBE]=8'h21; mem['h0EBF]=8'hD0;
    mem['h0EC0]=8'h0E; mem['h0EC1]=8'h3A; mem['h0EC2]=8'hF2; mem['h0EC3]=8'h80;
    mem['h0EC4]=8'h1F; mem['h0EC5]=8'h7A; mem['h0EC6]=8'h17; mem['h0EC7]=8'h5F;
    mem['h0EC8]=8'h16; mem['h0EC9]=8'h64; mem['h0ECA]=8'h78; mem['h0ECB]=8'hBA;
    mem['h0ECC]=8'hD0; mem['h0ECD]=8'hC3; mem['h0ECE]=8'hBF; mem['h0ECF]=8'h0D;
    mem['h0ED0]=8'hD2; mem['h0ED1]=8'h0E; mem['h0ED2]=8'h79; mem['h0ED3]=8'hB7;
    mem['h0ED4]=8'h1F; mem['h0ED5]=8'hC1; mem['h0ED6]=8'hD1; mem['h0ED7]=8'hF5;
    mem['h0ED8]=8'hCD; mem['h0ED9]=8'h52; mem['h0EDA]=8'h0D; mem['h0EDB]=8'h21;
    mem['h0EDC]=8'h14; mem['h0EDD]=8'h0F; mem['h0EDE]=8'hE5; mem['h0EDF]=8'hCA;
    mem['h0EE0]=8'hAA; mem['h0EE1]=8'h17; mem['h0EE2]=8'hAF; mem['h0EE3]=8'h32;
    mem['h0EE4]=8'hF2; mem['h0EE5]=8'h80; mem['h0EE6]=8'hD5; mem['h0EE7]=8'hCD;
    mem['h0EE8]=8'h69; mem['h0EE9]=8'h13; mem['h0EEA]=8'h7E; mem['h0EEB]=8'h23;
    mem['h0EEC]=8'h23; mem['h0EED]=8'h4E; mem['h0EEE]=8'h23; mem['h0EEF]=8'h46;
    mem['h0EF0]=8'hD1; mem['h0EF1]=8'hC5; mem['h0EF2]=8'hF5; mem['h0EF3]=8'hCD;
    mem['h0EF4]=8'h6D; mem['h0EF5]=8'h13; mem['h0EF6]=8'hCD; mem['h0EF7]=8'h7E;
    mem['h0EF8]=8'h17; mem['h0EF9]=8'hF1; mem['h0EFA]=8'h57; mem['h0EFB]=8'hE1;
    mem['h0EFC]=8'h7B; mem['h0EFD]=8'hB2; mem['h0EFE]=8'hC8; mem['h0EFF]=8'h7A;
    mem['h0F00]=8'hD6; mem['h0F01]=8'h01; mem['h0F02]=8'hD8; mem['h0F03]=8'hAF;
    mem['h0F04]=8'hBB; mem['h0F05]=8'h3C; mem['h0F06]=8'hD0; mem['h0F07]=8'h15;
    mem['h0F08]=8'h1D; mem['h0F09]=8'h0A; mem['h0F0A]=8'hBE; mem['h0F0B]=8'h23;
    mem['h0F0C]=8'h03; mem['h0F0D]=8'hCA; mem['h0F0E]=8'hFC; mem['h0F0F]=8'h0E;
    mem['h0F10]=8'h3F; mem['h0F11]=8'hC3; mem['h0F12]=8'h3A; mem['h0F13]=8'h17;
    mem['h0F14]=8'h3C; mem['h0F15]=8'h8F; mem['h0F16]=8'hC1; mem['h0F17]=8'hA0;
    mem['h0F18]=8'hC6; mem['h0F19]=8'hFF; mem['h0F1A]=8'h9F; mem['h0F1B]=8'hC3;
    mem['h0F1C]=8'h41; mem['h0F1D]=8'h17; mem['h0F1E]=8'h16; mem['h0F1F]=8'h5A;
    mem['h0F20]=8'hCD; mem['h0F21]=8'h62; mem['h0F22]=8'h0D; mem['h0F23]=8'hCD;
    mem['h0F24]=8'h50; mem['h0F25]=8'h0D; mem['h0F26]=8'hCD; mem['h0F27]=8'h92;
    mem['h0F28]=8'h09; mem['h0F29]=8'h7B; mem['h0F2A]=8'h2F; mem['h0F2B]=8'h4F;
    mem['h0F2C]=8'h7A; mem['h0F2D]=8'h2F; mem['h0F2E]=8'hCD; mem['h0F2F]=8'h07;
    mem['h0F30]=8'h11; mem['h0F31]=8'hC1; mem['h0F32]=8'hC3; mem['h0F33]=8'h6E;
    mem['h0F34]=8'h0D; mem['h0F35]=8'h2B; mem['h0F36]=8'hCD; mem['h0F37]=8'hE0;
    mem['h0F38]=8'h08; mem['h0F39]=8'hC8; mem['h0F3A]=8'hCD; mem['h0F3B]=8'h56;
    mem['h0F3C]=8'h07; mem['h0F3D]=8'h2C; mem['h0F3E]=8'h01; mem['h0F3F]=8'h35;
    mem['h0F40]=8'h0F; mem['h0F41]=8'hC5; mem['h0F42]=8'hF6; mem['h0F43]=8'hAF;
    mem['h0F44]=8'h32; mem['h0F45]=8'hF1; mem['h0F46]=8'h80; mem['h0F47]=8'h46;
    mem['h0F48]=8'hCD; mem['h0F49]=8'h7E; mem['h0F4A]=8'h09; mem['h0F4B]=8'hDA;
    mem['h0F4C]=8'h88; mem['h0F4D]=8'h04; mem['h0F4E]=8'hAF; mem['h0F4F]=8'h4F;
    mem['h0F50]=8'h32; mem['h0F51]=8'hF2; mem['h0F52]=8'h80; mem['h0F53]=8'hCD;
    mem['h0F54]=8'hE0; mem['h0F55]=8'h08; mem['h0F56]=8'hDA; mem['h0F57]=8'h5F;
    mem['h0F58]=8'h0F; mem['h0F59]=8'hCD; mem['h0F5A]=8'h7E; mem['h0F5B]=8'h09;
    mem['h0F5C]=8'hDA; mem['h0F5D]=8'h6C; mem['h0F5E]=8'h0F; mem['h0F5F]=8'h4F;
    mem['h0F60]=8'hCD; mem['h0F61]=8'hE0; mem['h0F62]=8'h08; mem['h0F63]=8'hDA;
    mem['h0F64]=8'h60; mem['h0F65]=8'h0F; mem['h0F66]=8'hCD; mem['h0F67]=8'h7E;
    mem['h0F68]=8'h09; mem['h0F69]=8'hD2; mem['h0F6A]=8'h60; mem['h0F6B]=8'h0F;
    mem['h0F6C]=8'hD6; mem['h0F6D]=8'h24; mem['h0F6E]=8'hC2; mem['h0F6F]=8'h7B;
    mem['h0F70]=8'h0F; mem['h0F71]=8'h3C; mem['h0F72]=8'h32; mem['h0F73]=8'hF2;
    mem['h0F74]=8'h80; mem['h0F75]=8'h0F; mem['h0F76]=8'h81; mem['h0F77]=8'h4F;
    mem['h0F78]=8'hCD; mem['h0F79]=8'hE0; mem['h0F7A]=8'h08; mem['h0F7B]=8'h3A;
    mem['h0F7C]=8'h10; mem['h0F7D]=8'h81; mem['h0F7E]=8'h3D; mem['h0F7F]=8'hCA;
    mem['h0F80]=8'h28; mem['h0F81]=8'h10; mem['h0F82]=8'hF2; mem['h0F83]=8'h8B;
    mem['h0F84]=8'h0F; mem['h0F85]=8'h7E; mem['h0F86]=8'hD6; mem['h0F87]=8'h28;
    mem['h0F88]=8'hCA; mem['h0F89]=8'h00; mem['h0F8A]=8'h10; mem['h0F8B]=8'hAF;
    mem['h0F8C]=8'h32; mem['h0F8D]=8'h10; mem['h0F8E]=8'h81; mem['h0F8F]=8'hE5;
    mem['h0F90]=8'h50; mem['h0F91]=8'h59; mem['h0F92]=8'h2A; mem['h0F93]=8'h23;
    mem['h0F94]=8'h81; mem['h0F95]=8'hCD; mem['h0F96]=8'h50; mem['h0F97]=8'h07;
    mem['h0F98]=8'h11; mem['h0F99]=8'h25; mem['h0F9A]=8'h81; mem['h0F9B]=8'hCA;
    mem['h0F9C]=8'h70; mem['h0F9D]=8'h16; mem['h0F9E]=8'h2A; mem['h0F9F]=8'h1D;
    mem['h0FA0]=8'h81; mem['h0FA1]=8'hEB; mem['h0FA2]=8'h2A; mem['h0FA3]=8'h1B;
    mem['h0FA4]=8'h81; mem['h0FA5]=8'hCD; mem['h0FA6]=8'h50; mem['h0FA7]=8'h07;
    mem['h0FA8]=8'hCA; mem['h0FA9]=8'hBE; mem['h0FAA]=8'h0F; mem['h0FAB]=8'h79;
    mem['h0FAC]=8'h96; mem['h0FAD]=8'h23; mem['h0FAE]=8'hC2; mem['h0FAF]=8'hB3;
    mem['h0FB0]=8'h0F; mem['h0FB1]=8'h78; mem['h0FB2]=8'h96; mem['h0FB3]=8'h23;
    mem['h0FB4]=8'hCA; mem['h0FB5]=8'hF2; mem['h0FB6]=8'h0F; mem['h0FB7]=8'h23;
    mem['h0FB8]=8'h23; mem['h0FB9]=8'h23; mem['h0FBA]=8'h23; mem['h0FBB]=8'hC3;
    mem['h0FBC]=8'hA5; mem['h0FBD]=8'h0F; mem['h0FBE]=8'hE1; mem['h0FBF]=8'hE3;
    mem['h0FC0]=8'hD5; mem['h0FC1]=8'h11; mem['h0FC2]=8'h40; mem['h0FC3]=8'h0E;
    mem['h0FC4]=8'hCD; mem['h0FC5]=8'h50; mem['h0FC6]=8'h07; mem['h0FC7]=8'hD1;
    mem['h0FC8]=8'hCA; mem['h0FC9]=8'hF5; mem['h0FCA]=8'h0F; mem['h0FCB]=8'hE3;
    mem['h0FCC]=8'hE5; mem['h0FCD]=8'hC5; mem['h0FCE]=8'h01; mem['h0FCF]=8'h06;
    mem['h0FD0]=8'h00; mem['h0FD1]=8'h2A; mem['h0FD2]=8'h1F; mem['h0FD3]=8'h81;
    mem['h0FD4]=8'hE5; mem['h0FD5]=8'h09; mem['h0FD6]=8'hC1; mem['h0FD7]=8'hE5;
    mem['h0FD8]=8'hCD; mem['h0FD9]=8'h54; mem['h0FDA]=8'h04; mem['h0FDB]=8'hE1;
    mem['h0FDC]=8'h22; mem['h0FDD]=8'h1F; mem['h0FDE]=8'h81; mem['h0FDF]=8'h60;
    mem['h0FE0]=8'h69; mem['h0FE1]=8'h22; mem['h0FE2]=8'h1D; mem['h0FE3]=8'h81;
    mem['h0FE4]=8'h2B; mem['h0FE5]=8'h36; mem['h0FE6]=8'h00; mem['h0FE7]=8'hCD;
    mem['h0FE8]=8'h50; mem['h0FE9]=8'h07; mem['h0FEA]=8'hC2; mem['h0FEB]=8'hE4;
    mem['h0FEC]=8'h0F; mem['h0FED]=8'hD1; mem['h0FEE]=8'h73; mem['h0FEF]=8'h23;
    mem['h0FF0]=8'h72; mem['h0FF1]=8'h23; mem['h0FF2]=8'hEB; mem['h0FF3]=8'hE1;
    mem['h0FF4]=8'hC9; mem['h0FF5]=8'h32; mem['h0FF6]=8'h2C; mem['h0FF7]=8'h81;
    mem['h0FF8]=8'h21; mem['h0FF9]=8'h24; mem['h0FFA]=8'h04; mem['h0FFB]=8'h22;
    mem['h0FFC]=8'h29; mem['h0FFD]=8'h81; mem['h0FFE]=8'hE1; mem['h0FFF]=8'hC9;
    mem['h1000]=8'hE5; mem['h1001]=8'h2A; mem['h1002]=8'hF1; mem['h1003]=8'h80;
    mem['h1004]=8'hE3; mem['h1005]=8'h57; mem['h1006]=8'hD5; mem['h1007]=8'hC5;
    mem['h1008]=8'hCD; mem['h1009]=8'h86; mem['h100A]=8'h09; mem['h100B]=8'hC1;
    mem['h100C]=8'hF1; mem['h100D]=8'hEB; mem['h100E]=8'hE3; mem['h100F]=8'hE5;
    mem['h1010]=8'hEB; mem['h1011]=8'h3C; mem['h1012]=8'h57; mem['h1013]=8'h7E;
    mem['h1014]=8'hFE; mem['h1015]=8'h2C; mem['h1016]=8'hCA; mem['h1017]=8'h06;
    mem['h1018]=8'h10; mem['h1019]=8'hCD; mem['h101A]=8'h56; mem['h101B]=8'h07;
    mem['h101C]=8'h29; mem['h101D]=8'h22; mem['h101E]=8'h15; mem['h101F]=8'h81;
    mem['h1020]=8'hE1; mem['h1021]=8'h22; mem['h1022]=8'hF1; mem['h1023]=8'h80;
    mem['h1024]=8'h1E; mem['h1025]=8'h00; mem['h1026]=8'hD5; mem['h1027]=8'h11;
    mem['h1028]=8'hE5; mem['h1029]=8'hF5; mem['h102A]=8'h2A; mem['h102B]=8'h1D;
    mem['h102C]=8'h81; mem['h102D]=8'h3E; mem['h102E]=8'h19; mem['h102F]=8'hEB;
    mem['h1030]=8'h2A; mem['h1031]=8'h1F; mem['h1032]=8'h81; mem['h1033]=8'hEB;
    mem['h1034]=8'hCD; mem['h1035]=8'h50; mem['h1036]=8'h07; mem['h1037]=8'hCA;
    mem['h1038]=8'h60; mem['h1039]=8'h10; mem['h103A]=8'h7E; mem['h103B]=8'hB9;
    mem['h103C]=8'h23; mem['h103D]=8'hC2; mem['h103E]=8'h42; mem['h103F]=8'h10;
    mem['h1040]=8'h7E; mem['h1041]=8'hB8; mem['h1042]=8'h23; mem['h1043]=8'h5E;
    mem['h1044]=8'h23; mem['h1045]=8'h56; mem['h1046]=8'h23; mem['h1047]=8'hC2;
    mem['h1048]=8'h2E; mem['h1049]=8'h10; mem['h104A]=8'h3A; mem['h104B]=8'hF1;
    mem['h104C]=8'h80; mem['h104D]=8'hB7; mem['h104E]=8'hC2; mem['h104F]=8'h91;
    mem['h1050]=8'h04; mem['h1051]=8'hF1; mem['h1052]=8'h44; mem['h1053]=8'h4D;
    mem['h1054]=8'hCA; mem['h1055]=8'h70; mem['h1056]=8'h16; mem['h1057]=8'h96;
    mem['h1058]=8'hCA; mem['h1059]=8'hBE; mem['h105A]=8'h10; mem['h105B]=8'h1E;
    mem['h105C]=8'h10; mem['h105D]=8'hC3; mem['h105E]=8'h9C; mem['h105F]=8'h04;
    mem['h1060]=8'h11; mem['h1061]=8'h04; mem['h1062]=8'h00; mem['h1063]=8'hF1;
    mem['h1064]=8'hCA; mem['h1065]=8'hA7; mem['h1066]=8'h09; mem['h1067]=8'h71;
    mem['h1068]=8'h23; mem['h1069]=8'h70; mem['h106A]=8'h23; mem['h106B]=8'h4F;
    mem['h106C]=8'hCD; mem['h106D]=8'h65; mem['h106E]=8'h04; mem['h106F]=8'h23;
    mem['h1070]=8'h23; mem['h1071]=8'h22; mem['h1072]=8'h0A; mem['h1073]=8'h81;
    mem['h1074]=8'h71; mem['h1075]=8'h23; mem['h1076]=8'h3A; mem['h1077]=8'hF1;
    mem['h1078]=8'h80; mem['h1079]=8'h17; mem['h107A]=8'h79; mem['h107B]=8'h01;
    mem['h107C]=8'h0B; mem['h107D]=8'h00; mem['h107E]=8'hD2; mem['h107F]=8'h83;
    mem['h1080]=8'h10; mem['h1081]=8'hC1; mem['h1082]=8'h03; mem['h1083]=8'h71;
    mem['h1084]=8'h23; mem['h1085]=8'h70; mem['h1086]=8'h23; mem['h1087]=8'hF5;
    mem['h1088]=8'hE5; mem['h1089]=8'hCD; mem['h108A]=8'h1B; mem['h108B]=8'h18;
    mem['h108C]=8'hEB; mem['h108D]=8'hE1; mem['h108E]=8'hF1; mem['h108F]=8'h3D;
    mem['h1090]=8'hC2; mem['h1091]=8'h7B; mem['h1092]=8'h10; mem['h1093]=8'hF5;
    mem['h1094]=8'h42; mem['h1095]=8'h4B; mem['h1096]=8'hEB; mem['h1097]=8'h19;
    mem['h1098]=8'hDA; mem['h1099]=8'h7D; mem['h109A]=8'h04; mem['h109B]=8'hCD;
    mem['h109C]=8'h6E; mem['h109D]=8'h04; mem['h109E]=8'h22; mem['h109F]=8'h1F;
    mem['h10A0]=8'h81; mem['h10A1]=8'h2B; mem['h10A2]=8'h36; mem['h10A3]=8'h00;
    mem['h10A4]=8'hCD; mem['h10A5]=8'h50; mem['h10A6]=8'h07; mem['h10A7]=8'hC2;
    mem['h10A8]=8'hA1; mem['h10A9]=8'h10; mem['h10AA]=8'h03; mem['h10AB]=8'h57;
    mem['h10AC]=8'h2A; mem['h10AD]=8'h0A; mem['h10AE]=8'h81; mem['h10AF]=8'h5E;
    mem['h10B0]=8'hEB; mem['h10B1]=8'h29; mem['h10B2]=8'h09; mem['h10B3]=8'hEB;
    mem['h10B4]=8'h2B; mem['h10B5]=8'h2B; mem['h10B6]=8'h73; mem['h10B7]=8'h23;
    mem['h10B8]=8'h72; mem['h10B9]=8'h23; mem['h10BA]=8'hF1; mem['h10BB]=8'hDA;
    mem['h10BC]=8'hE2; mem['h10BD]=8'h10; mem['h10BE]=8'h47; mem['h10BF]=8'h4F;
    mem['h10C0]=8'h7E; mem['h10C1]=8'h23; mem['h10C2]=8'h16; mem['h10C3]=8'hE1;
    mem['h10C4]=8'h5E; mem['h10C5]=8'h23; mem['h10C6]=8'h56; mem['h10C7]=8'h23;
    mem['h10C8]=8'hE3; mem['h10C9]=8'hF5; mem['h10CA]=8'hCD; mem['h10CB]=8'h50;
    mem['h10CC]=8'h07; mem['h10CD]=8'hD2; mem['h10CE]=8'h5B; mem['h10CF]=8'h10;
    mem['h10D0]=8'hE5; mem['h10D1]=8'hCD; mem['h10D2]=8'h1B; mem['h10D3]=8'h18;
    mem['h10D4]=8'hD1; mem['h10D5]=8'h19; mem['h10D6]=8'hF1; mem['h10D7]=8'h3D;
    mem['h10D8]=8'h44; mem['h10D9]=8'h4D; mem['h10DA]=8'hC2; mem['h10DB]=8'hC3;
    mem['h10DC]=8'h10; mem['h10DD]=8'h29; mem['h10DE]=8'h29; mem['h10DF]=8'hC1;
    mem['h10E0]=8'h09; mem['h10E1]=8'hEB; mem['h10E2]=8'h2A; mem['h10E3]=8'h15;
    mem['h10E4]=8'h81; mem['h10E5]=8'hC9; mem['h10E6]=8'h2A; mem['h10E7]=8'h1F;
    mem['h10E8]=8'h81; mem['h10E9]=8'hEB; mem['h10EA]=8'h21; mem['h10EB]=8'h00;
    mem['h10EC]=8'h00; mem['h10ED]=8'h39; mem['h10EE]=8'h3A; mem['h10EF]=8'hF2;
    mem['h10F0]=8'h80; mem['h10F1]=8'hB7; mem['h10F2]=8'hCA; mem['h10F3]=8'h02;
    mem['h10F4]=8'h11; mem['h10F5]=8'hCD; mem['h10F6]=8'h69; mem['h10F7]=8'h13;
    mem['h10F8]=8'hCD; mem['h10F9]=8'h69; mem['h10FA]=8'h12; mem['h10FB]=8'h2A;
    mem['h10FC]=8'h9F; mem['h10FD]=8'h80; mem['h10FE]=8'hEB; mem['h10FF]=8'h2A;
    mem['h1100]=8'h08; mem['h1101]=8'h81; mem['h1102]=8'h7D; mem['h1103]=8'h93;
    mem['h1104]=8'h4F; mem['h1105]=8'h7C; mem['h1106]=8'h9A; mem['h1107]=8'h41;
    mem['h1108]=8'h50; mem['h1109]=8'h1E; mem['h110A]=8'h00; mem['h110B]=8'h21;
    mem['h110C]=8'hF2; mem['h110D]=8'h80; mem['h110E]=8'h73; mem['h110F]=8'h06;
    mem['h1110]=8'h90; mem['h1111]=8'hC3; mem['h1112]=8'h46; mem['h1113]=8'h17;
    mem['h1114]=8'h3A; mem['h1115]=8'hF0; mem['h1116]=8'h80; mem['h1117]=8'h47;
    mem['h1118]=8'hAF; mem['h1119]=8'hC3; mem['h111A]=8'h08; mem['h111B]=8'h11;
    mem['h111C]=8'hCD; mem['h111D]=8'h9F; mem['h111E]=8'h11; mem['h111F]=8'hCD;
    mem['h1120]=8'h91; mem['h1121]=8'h11; mem['h1122]=8'h01; mem['h1123]=8'h77;
    mem['h1124]=8'h0A; mem['h1125]=8'hC5; mem['h1126]=8'hD5; mem['h1127]=8'hCD;
    mem['h1128]=8'h56; mem['h1129]=8'h07; mem['h112A]=8'h28; mem['h112B]=8'hCD;
    mem['h112C]=8'h43; mem['h112D]=8'h0F; mem['h112E]=8'hE5; mem['h112F]=8'hEB;
    mem['h1130]=8'h2B; mem['h1131]=8'h56; mem['h1132]=8'h2B; mem['h1133]=8'h5E;
    mem['h1134]=8'hE1; mem['h1135]=8'hCD; mem['h1136]=8'h50; mem['h1137]=8'h0D;
    mem['h1138]=8'hCD; mem['h1139]=8'h56; mem['h113A]=8'h07; mem['h113B]=8'h29;
    mem['h113C]=8'hCD; mem['h113D]=8'h56; mem['h113E]=8'h07; mem['h113F]=8'hB4;
    mem['h1140]=8'h44; mem['h1141]=8'h4D; mem['h1142]=8'hE3; mem['h1143]=8'h71;
    mem['h1144]=8'h23; mem['h1145]=8'h70; mem['h1146]=8'hC3; mem['h1147]=8'hDE;
    mem['h1148]=8'h11; mem['h1149]=8'hCD; mem['h114A]=8'h9F; mem['h114B]=8'h11;
    mem['h114C]=8'hD5; mem['h114D]=8'hCD; mem['h114E]=8'h24; mem['h114F]=8'h0E;
    mem['h1150]=8'hCD; mem['h1151]=8'h50; mem['h1152]=8'h0D; mem['h1153]=8'hE3;
    mem['h1154]=8'h5E; mem['h1155]=8'h23; mem['h1156]=8'h56; mem['h1157]=8'h23;
    mem['h1158]=8'h7A; mem['h1159]=8'hB3; mem['h115A]=8'hCA; mem['h115B]=8'h94;
    mem['h115C]=8'h04; mem['h115D]=8'h7E; mem['h115E]=8'h23; mem['h115F]=8'h66;
    mem['h1160]=8'h6F; mem['h1161]=8'hE5; mem['h1162]=8'h2A; mem['h1163]=8'h23;
    mem['h1164]=8'h81; mem['h1165]=8'hE3; mem['h1166]=8'h22; mem['h1167]=8'h23;
    mem['h1168]=8'h81; mem['h1169]=8'h2A; mem['h116A]=8'h27; mem['h116B]=8'h81;
    mem['h116C]=8'hE5; mem['h116D]=8'h2A; mem['h116E]=8'h25; mem['h116F]=8'h81;
    mem['h1170]=8'hE5; mem['h1171]=8'h21; mem['h1172]=8'h25; mem['h1173]=8'h81;
    mem['h1174]=8'hD5; mem['h1175]=8'hCD; mem['h1176]=8'h87; mem['h1177]=8'h17;
    mem['h1178]=8'hE1; mem['h1179]=8'hCD; mem['h117A]=8'h4D; mem['h117B]=8'h0D;
    mem['h117C]=8'h2B; mem['h117D]=8'hCD; mem['h117E]=8'hE0; mem['h117F]=8'h08;
    mem['h1180]=8'hC2; mem['h1181]=8'h88; mem['h1182]=8'h04; mem['h1183]=8'hE1;
    mem['h1184]=8'h22; mem['h1185]=8'h25; mem['h1186]=8'h81; mem['h1187]=8'hE1;
    mem['h1188]=8'h22; mem['h1189]=8'h27; mem['h118A]=8'h81; mem['h118B]=8'hE1;
    mem['h118C]=8'h22; mem['h118D]=8'h23; mem['h118E]=8'h81; mem['h118F]=8'hE1;
    mem['h1190]=8'hC9; mem['h1191]=8'hE5; mem['h1192]=8'h2A; mem['h1193]=8'hA1;
    mem['h1194]=8'h80; mem['h1195]=8'h23; mem['h1196]=8'h7C; mem['h1197]=8'hB5;
    mem['h1198]=8'hE1; mem['h1199]=8'hC0; mem['h119A]=8'h1E; mem['h119B]=8'h16;
    mem['h119C]=8'hC3; mem['h119D]=8'h9C; mem['h119E]=8'h04; mem['h119F]=8'hCD;
    mem['h11A0]=8'h56; mem['h11A1]=8'h07; mem['h11A2]=8'hA7; mem['h11A3]=8'h3E;
    mem['h11A4]=8'h80; mem['h11A5]=8'h32; mem['h11A6]=8'h10; mem['h11A7]=8'h81;
    mem['h11A8]=8'hB6; mem['h11A9]=8'h47; mem['h11AA]=8'hCD; mem['h11AB]=8'h48;
    mem['h11AC]=8'h0F; mem['h11AD]=8'hC3; mem['h11AE]=8'h50; mem['h11AF]=8'h0D;
    mem['h11B0]=8'hCD; mem['h11B1]=8'h50; mem['h11B2]=8'h0D; mem['h11B3]=8'hCD;
    mem['h11B4]=8'hD4; mem['h11B5]=8'h18; mem['h11B6]=8'hCD; mem['h11B7]=8'hE4;
    mem['h11B8]=8'h11; mem['h11B9]=8'hCD; mem['h11BA]=8'h69; mem['h11BB]=8'h13;
    mem['h11BC]=8'h01; mem['h11BD]=8'hC4; mem['h11BE]=8'h13; mem['h11BF]=8'hC5;
    mem['h11C0]=8'h7E; mem['h11C1]=8'h23; mem['h11C2]=8'h23; mem['h11C3]=8'hE5;
    mem['h11C4]=8'hCD; mem['h11C5]=8'h3F; mem['h11C6]=8'h12; mem['h11C7]=8'hE1;
    mem['h11C8]=8'h4E; mem['h11C9]=8'h23; mem['h11CA]=8'h46; mem['h11CB]=8'hCD;
    mem['h11CC]=8'hD8; mem['h11CD]=8'h11; mem['h11CE]=8'hE5; mem['h11CF]=8'h6F;
    mem['h11D0]=8'hCD; mem['h11D1]=8'h5C; mem['h11D2]=8'h13; mem['h11D3]=8'hD1;
    mem['h11D4]=8'hC9; mem['h11D5]=8'hCD; mem['h11D6]=8'h3F; mem['h11D7]=8'h12;
    mem['h11D8]=8'h21; mem['h11D9]=8'h04; mem['h11DA]=8'h81; mem['h11DB]=8'hE5;
    mem['h11DC]=8'h77; mem['h11DD]=8'h23; mem['h11DE]=8'h23; mem['h11DF]=8'h73;
    mem['h11E0]=8'h23; mem['h11E1]=8'h72; mem['h11E2]=8'hE1; mem['h11E3]=8'hC9;
    mem['h11E4]=8'h2B; mem['h11E5]=8'h06; mem['h11E6]=8'h22; mem['h11E7]=8'h50;
    mem['h11E8]=8'hE5; mem['h11E9]=8'h0E; mem['h11EA]=8'hFF; mem['h11EB]=8'h23;
    mem['h11EC]=8'h7E; mem['h11ED]=8'h0C; mem['h11EE]=8'hB7; mem['h11EF]=8'hCA;
    mem['h11F0]=8'hFA; mem['h11F1]=8'h11; mem['h11F2]=8'hBA; mem['h11F3]=8'hCA;
    mem['h11F4]=8'hFA; mem['h11F5]=8'h11; mem['h11F6]=8'hB8; mem['h11F7]=8'hC2;
    mem['h11F8]=8'hEB; mem['h11F9]=8'h11; mem['h11FA]=8'hFE; mem['h11FB]=8'h22;
    mem['h11FC]=8'hCC; mem['h11FD]=8'hE0; mem['h11FE]=8'h08; mem['h11FF]=8'hE3;
    mem['h1200]=8'h23; mem['h1201]=8'hEB; mem['h1202]=8'h79; mem['h1203]=8'hCD;
    mem['h1204]=8'hD8; mem['h1205]=8'h11; mem['h1206]=8'h11; mem['h1207]=8'h04;
    mem['h1208]=8'h81; mem['h1209]=8'h2A; mem['h120A]=8'hF6; mem['h120B]=8'h80;
    mem['h120C]=8'h22; mem['h120D]=8'h29; mem['h120E]=8'h81; mem['h120F]=8'h3E;
    mem['h1210]=8'h01; mem['h1211]=8'h32; mem['h1212]=8'hF2; mem['h1213]=8'h80;
    mem['h1214]=8'hCD; mem['h1215]=8'h8A; mem['h1216]=8'h17; mem['h1217]=8'hCD;
    mem['h1218]=8'h50; mem['h1219]=8'h07; mem['h121A]=8'h22; mem['h121B]=8'hF6;
    mem['h121C]=8'h80; mem['h121D]=8'hE1; mem['h121E]=8'h7E; mem['h121F]=8'hC0;
    mem['h1220]=8'h1E; mem['h1221]=8'h1E; mem['h1222]=8'hC3; mem['h1223]=8'h9C;
    mem['h1224]=8'h04; mem['h1225]=8'h23; mem['h1226]=8'hCD; mem['h1227]=8'hE4;
    mem['h1228]=8'h11; mem['h1229]=8'hCD; mem['h122A]=8'h69; mem['h122B]=8'h13;
    mem['h122C]=8'hCD; mem['h122D]=8'h7E; mem['h122E]=8'h17; mem['h122F]=8'h1C;
    mem['h1230]=8'h1D; mem['h1231]=8'hC8; mem['h1232]=8'h0A; mem['h1233]=8'hCD;
    mem['h1234]=8'h61; mem['h1235]=8'h07; mem['h1236]=8'hFE; mem['h1237]=8'h0D;
    mem['h1238]=8'hCC; mem['h1239]=8'h92; mem['h123A]=8'h0B; mem['h123B]=8'h03;
    mem['h123C]=8'hC3; mem['h123D]=8'h30; mem['h123E]=8'h12; mem['h123F]=8'hB7;
    mem['h1240]=8'h0E; mem['h1241]=8'hF1; mem['h1242]=8'hF5; mem['h1243]=8'h2A;
    mem['h1244]=8'h9F; mem['h1245]=8'h80; mem['h1246]=8'hEB; mem['h1247]=8'h2A;
    mem['h1248]=8'h08; mem['h1249]=8'h81; mem['h124A]=8'h2F; mem['h124B]=8'h4F;
    mem['h124C]=8'h06; mem['h124D]=8'hFF; mem['h124E]=8'h09; mem['h124F]=8'h23;
    mem['h1250]=8'hCD; mem['h1251]=8'h50; mem['h1252]=8'h07; mem['h1253]=8'hDA;
    mem['h1254]=8'h5D; mem['h1255]=8'h12; mem['h1256]=8'h22; mem['h1257]=8'h08;
    mem['h1258]=8'h81; mem['h1259]=8'h23; mem['h125A]=8'hEB; mem['h125B]=8'hF1;
    mem['h125C]=8'hC9; mem['h125D]=8'hF1; mem['h125E]=8'h1E; mem['h125F]=8'h1A;
    mem['h1260]=8'hCA; mem['h1261]=8'h9C; mem['h1262]=8'h04; mem['h1263]=8'hBF;
    mem['h1264]=8'hF5; mem['h1265]=8'h01; mem['h1266]=8'h41; mem['h1267]=8'h12;
    mem['h1268]=8'hC5; mem['h1269]=8'h2A; mem['h126A]=8'hF4; mem['h126B]=8'h80;
    mem['h126C]=8'h22; mem['h126D]=8'h08; mem['h126E]=8'h81; mem['h126F]=8'h21;
    mem['h1270]=8'h00; mem['h1271]=8'h00; mem['h1272]=8'hE5; mem['h1273]=8'h2A;
    mem['h1274]=8'h9F; mem['h1275]=8'h80; mem['h1276]=8'hE5; mem['h1277]=8'h21;
    mem['h1278]=8'hF8; mem['h1279]=8'h80; mem['h127A]=8'hEB; mem['h127B]=8'h2A;
    mem['h127C]=8'hF6; mem['h127D]=8'h80; mem['h127E]=8'hEB; mem['h127F]=8'hCD;
    mem['h1280]=8'h50; mem['h1281]=8'h07; mem['h1282]=8'h01; mem['h1283]=8'h7A;
    mem['h1284]=8'h12; mem['h1285]=8'hC2; mem['h1286]=8'hCE; mem['h1287]=8'h12;
    mem['h1288]=8'h2A; mem['h1289]=8'h1B; mem['h128A]=8'h81; mem['h128B]=8'hEB;
    mem['h128C]=8'h2A; mem['h128D]=8'h1D; mem['h128E]=8'h81; mem['h128F]=8'hEB;
    mem['h1290]=8'hCD; mem['h1291]=8'h50; mem['h1292]=8'h07; mem['h1293]=8'hCA;
    mem['h1294]=8'hA1; mem['h1295]=8'h12; mem['h1296]=8'h7E; mem['h1297]=8'h23;
    mem['h1298]=8'h23; mem['h1299]=8'hB7; mem['h129A]=8'hCD; mem['h129B]=8'hD1;
    mem['h129C]=8'h12; mem['h129D]=8'hC3; mem['h129E]=8'h8B; mem['h129F]=8'h12;
    mem['h12A0]=8'hC1; mem['h12A1]=8'hEB; mem['h12A2]=8'h2A; mem['h12A3]=8'h1F;
    mem['h12A4]=8'h81; mem['h12A5]=8'hEB; mem['h12A6]=8'hCD; mem['h12A7]=8'h50;
    mem['h12A8]=8'h07; mem['h12A9]=8'hCA; mem['h12AA]=8'hF7; mem['h12AB]=8'h12;
    mem['h12AC]=8'hCD; mem['h12AD]=8'h7E; mem['h12AE]=8'h17; mem['h12AF]=8'h7B;
    mem['h12B0]=8'hE5; mem['h12B1]=8'h09; mem['h12B2]=8'hB7; mem['h12B3]=8'hF2;
    mem['h12B4]=8'hA0; mem['h12B5]=8'h12; mem['h12B6]=8'h22; mem['h12B7]=8'h0A;
    mem['h12B8]=8'h81; mem['h12B9]=8'hE1; mem['h12BA]=8'h4E; mem['h12BB]=8'h06;
    mem['h12BC]=8'h00; mem['h12BD]=8'h09; mem['h12BE]=8'h09; mem['h12BF]=8'h23;
    mem['h12C0]=8'hEB; mem['h12C1]=8'h2A; mem['h12C2]=8'h0A; mem['h12C3]=8'h81;
    mem['h12C4]=8'hEB; mem['h12C5]=8'hCD; mem['h12C6]=8'h50; mem['h12C7]=8'h07;
    mem['h12C8]=8'hCA; mem['h12C9]=8'hA1; mem['h12CA]=8'h12; mem['h12CB]=8'h01;
    mem['h12CC]=8'hC0; mem['h12CD]=8'h12; mem['h12CE]=8'hC5; mem['h12CF]=8'hF6;
    mem['h12D0]=8'h80; mem['h12D1]=8'h7E; mem['h12D2]=8'h23; mem['h12D3]=8'h23;
    mem['h12D4]=8'h5E; mem['h12D5]=8'h23; mem['h12D6]=8'h56; mem['h12D7]=8'h23;
    mem['h12D8]=8'hF0; mem['h12D9]=8'hB7; mem['h12DA]=8'hC8; mem['h12DB]=8'h44;
    mem['h12DC]=8'h4D; mem['h12DD]=8'h2A; mem['h12DE]=8'h08; mem['h12DF]=8'h81;
    mem['h12E0]=8'hCD; mem['h12E1]=8'h50; mem['h12E2]=8'h07; mem['h12E3]=8'h60;
    mem['h12E4]=8'h69; mem['h12E5]=8'hD8; mem['h12E6]=8'hE1; mem['h12E7]=8'hE3;
    mem['h12E8]=8'hCD; mem['h12E9]=8'h50; mem['h12EA]=8'h07; mem['h12EB]=8'hE3;
    mem['h12EC]=8'hE5; mem['h12ED]=8'h60; mem['h12EE]=8'h69; mem['h12EF]=8'hD0;
    mem['h12F0]=8'hC1; mem['h12F1]=8'hF1; mem['h12F2]=8'hF1; mem['h12F3]=8'hE5;
    mem['h12F4]=8'hD5; mem['h12F5]=8'hC5; mem['h12F6]=8'hC9; mem['h12F7]=8'hD1;
    mem['h12F8]=8'hE1; mem['h12F9]=8'h7D; mem['h12FA]=8'hB4; mem['h12FB]=8'hC8;
    mem['h12FC]=8'h2B; mem['h12FD]=8'h46; mem['h12FE]=8'h2B; mem['h12FF]=8'h4E;
    mem['h1300]=8'hE5; mem['h1301]=8'h2B; mem['h1302]=8'h2B; mem['h1303]=8'h6E;
    mem['h1304]=8'h26; mem['h1305]=8'h00; mem['h1306]=8'h09; mem['h1307]=8'h50;
    mem['h1308]=8'h59; mem['h1309]=8'h2B; mem['h130A]=8'h44; mem['h130B]=8'h4D;
    mem['h130C]=8'h2A; mem['h130D]=8'h08; mem['h130E]=8'h81; mem['h130F]=8'hCD;
    mem['h1310]=8'h57; mem['h1311]=8'h04; mem['h1312]=8'hE1; mem['h1313]=8'h71;
    mem['h1314]=8'h23; mem['h1315]=8'h70; mem['h1316]=8'h69; mem['h1317]=8'h60;
    mem['h1318]=8'h2B; mem['h1319]=8'hC3; mem['h131A]=8'h6C; mem['h131B]=8'h12;
    mem['h131C]=8'hC5; mem['h131D]=8'hE5; mem['h131E]=8'h2A; mem['h131F]=8'h29;
    mem['h1320]=8'h81; mem['h1321]=8'hE3; mem['h1322]=8'hCD; mem['h1323]=8'hD6;
    mem['h1324]=8'h0D; mem['h1325]=8'hE3; mem['h1326]=8'hCD; mem['h1327]=8'h51;
    mem['h1328]=8'h0D; mem['h1329]=8'h7E; mem['h132A]=8'hE5; mem['h132B]=8'h2A;
    mem['h132C]=8'h29; mem['h132D]=8'h81; mem['h132E]=8'hE5; mem['h132F]=8'h86;
    mem['h1330]=8'h1E; mem['h1331]=8'h1C; mem['h1332]=8'hDA; mem['h1333]=8'h9C;
    mem['h1334]=8'h04; mem['h1335]=8'hCD; mem['h1336]=8'hD5; mem['h1337]=8'h11;
    mem['h1338]=8'hD1; mem['h1339]=8'hCD; mem['h133A]=8'h6D; mem['h133B]=8'h13;
    mem['h133C]=8'hE3; mem['h133D]=8'hCD; mem['h133E]=8'h6C; mem['h133F]=8'h13;
    mem['h1340]=8'hE5; mem['h1341]=8'h2A; mem['h1342]=8'h06; mem['h1343]=8'h81;
    mem['h1344]=8'hEB; mem['h1345]=8'hCD; mem['h1346]=8'h53; mem['h1347]=8'h13;
    mem['h1348]=8'hCD; mem['h1349]=8'h53; mem['h134A]=8'h13; mem['h134B]=8'h21;
    mem['h134C]=8'h6B; mem['h134D]=8'h0D; mem['h134E]=8'hE3; mem['h134F]=8'hE5;
    mem['h1350]=8'hC3; mem['h1351]=8'h06; mem['h1352]=8'h12; mem['h1353]=8'hE1;
    mem['h1354]=8'hE3; mem['h1355]=8'h7E; mem['h1356]=8'h23; mem['h1357]=8'h23;
    mem['h1358]=8'h4E; mem['h1359]=8'h23; mem['h135A]=8'h46; mem['h135B]=8'h6F;
    mem['h135C]=8'h2C; mem['h135D]=8'h2D; mem['h135E]=8'hC8; mem['h135F]=8'h0A;
    mem['h1360]=8'h12; mem['h1361]=8'h03; mem['h1362]=8'h13; mem['h1363]=8'hC3;
    mem['h1364]=8'h5D; mem['h1365]=8'h13; mem['h1366]=8'hCD; mem['h1367]=8'h51;
    mem['h1368]=8'h0D; mem['h1369]=8'h2A; mem['h136A]=8'h29; mem['h136B]=8'h81;
    mem['h136C]=8'hEB; mem['h136D]=8'hCD; mem['h136E]=8'h87; mem['h136F]=8'h13;
    mem['h1370]=8'hEB; mem['h1371]=8'hC0; mem['h1372]=8'hD5; mem['h1373]=8'h50;
    mem['h1374]=8'h59; mem['h1375]=8'h1B; mem['h1376]=8'h4E; mem['h1377]=8'h2A;
    mem['h1378]=8'h08; mem['h1379]=8'h81; mem['h137A]=8'hCD; mem['h137B]=8'h50;
    mem['h137C]=8'h07; mem['h137D]=8'hC2; mem['h137E]=8'h85; mem['h137F]=8'h13;
    mem['h1380]=8'h47; mem['h1381]=8'h09; mem['h1382]=8'h22; mem['h1383]=8'h08;
    mem['h1384]=8'h81; mem['h1385]=8'hE1; mem['h1386]=8'hC9; mem['h1387]=8'h2A;
    mem['h1388]=8'hF6; mem['h1389]=8'h80; mem['h138A]=8'h2B; mem['h138B]=8'h46;
    mem['h138C]=8'h2B; mem['h138D]=8'h4E; mem['h138E]=8'h2B; mem['h138F]=8'h2B;
    mem['h1390]=8'hCD; mem['h1391]=8'h50; mem['h1392]=8'h07; mem['h1393]=8'hC0;
    mem['h1394]=8'h22; mem['h1395]=8'hF6; mem['h1396]=8'h80; mem['h1397]=8'hC9;
    mem['h1398]=8'h01; mem['h1399]=8'h17; mem['h139A]=8'h11; mem['h139B]=8'hC5;
    mem['h139C]=8'hCD; mem['h139D]=8'h66; mem['h139E]=8'h13; mem['h139F]=8'hAF;
    mem['h13A0]=8'h57; mem['h13A1]=8'h32; mem['h13A2]=8'hF2; mem['h13A3]=8'h80;
    mem['h13A4]=8'h7E; mem['h13A5]=8'hB7; mem['h13A6]=8'hC9; mem['h13A7]=8'h01;
    mem['h13A8]=8'h17; mem['h13A9]=8'h11; mem['h13AA]=8'hC5; mem['h13AB]=8'hCD;
    mem['h13AC]=8'h9C; mem['h13AD]=8'h13; mem['h13AE]=8'hCA; mem['h13AF]=8'hA7;
    mem['h13B0]=8'h09; mem['h13B1]=8'h23; mem['h13B2]=8'h23; mem['h13B3]=8'h5E;
    mem['h13B4]=8'h23; mem['h13B5]=8'h56; mem['h13B6]=8'h1A; mem['h13B7]=8'hC9;
    mem['h13B8]=8'h3E; mem['h13B9]=8'h01; mem['h13BA]=8'hCD; mem['h13BB]=8'hD5;
    mem['h13BC]=8'h11; mem['h13BD]=8'hCD; mem['h13BE]=8'hB1; mem['h13BF]=8'h14;
    mem['h13C0]=8'h2A; mem['h13C1]=8'h06; mem['h13C2]=8'h81; mem['h13C3]=8'h73;
    mem['h13C4]=8'hC1; mem['h13C5]=8'hC3; mem['h13C6]=8'h06; mem['h13C7]=8'h12;
    mem['h13C8]=8'hCD; mem['h13C9]=8'h61; mem['h13CA]=8'h14; mem['h13CB]=8'hAF;
    mem['h13CC]=8'hE3; mem['h13CD]=8'h4F; mem['h13CE]=8'hE5; mem['h13CF]=8'h7E;
    mem['h13D0]=8'hB8; mem['h13D1]=8'hDA; mem['h13D2]=8'hD6; mem['h13D3]=8'h13;
    mem['h13D4]=8'h78; mem['h13D5]=8'h11; mem['h13D6]=8'h0E; mem['h13D7]=8'h00;
    mem['h13D8]=8'hC5; mem['h13D9]=8'hCD; mem['h13DA]=8'h3F; mem['h13DB]=8'h12;
    mem['h13DC]=8'hC1; mem['h13DD]=8'hE1; mem['h13DE]=8'hE5; mem['h13DF]=8'h23;
    mem['h13E0]=8'h23; mem['h13E1]=8'h46; mem['h13E2]=8'h23; mem['h13E3]=8'h66;
    mem['h13E4]=8'h68; mem['h13E5]=8'h06; mem['h13E6]=8'h00; mem['h13E7]=8'h09;
    mem['h13E8]=8'h44; mem['h13E9]=8'h4D; mem['h13EA]=8'hCD; mem['h13EB]=8'hD8;
    mem['h13EC]=8'h11; mem['h13ED]=8'h6F; mem['h13EE]=8'hCD; mem['h13EF]=8'h5C;
    mem['h13F0]=8'h13; mem['h13F1]=8'hD1; mem['h13F2]=8'hCD; mem['h13F3]=8'h6D;
    mem['h13F4]=8'h13; mem['h13F5]=8'hC3; mem['h13F6]=8'h06; mem['h13F7]=8'h12;
    mem['h13F8]=8'hCD; mem['h13F9]=8'h61; mem['h13FA]=8'h14; mem['h13FB]=8'hD1;
    mem['h13FC]=8'hD5; mem['h13FD]=8'h1A; mem['h13FE]=8'h90; mem['h13FF]=8'hC3;
    mem['h1400]=8'hCC; mem['h1401]=8'h13; mem['h1402]=8'hEB; mem['h1403]=8'h7E;
    mem['h1404]=8'hCD; mem['h1405]=8'h66; mem['h1406]=8'h14; mem['h1407]=8'h04;
    mem['h1408]=8'h05; mem['h1409]=8'hCA; mem['h140A]=8'hA7; mem['h140B]=8'h09;
    mem['h140C]=8'hC5; mem['h140D]=8'h1E; mem['h140E]=8'hFF; mem['h140F]=8'hFE;
    mem['h1410]=8'h29; mem['h1411]=8'hCA; mem['h1412]=8'h1B; mem['h1413]=8'h14;
    mem['h1414]=8'hCD; mem['h1415]=8'h56; mem['h1416]=8'h07; mem['h1417]=8'h2C;
    mem['h1418]=8'hCD; mem['h1419]=8'hAE; mem['h141A]=8'h14; mem['h141B]=8'hCD;
    mem['h141C]=8'h56; mem['h141D]=8'h07; mem['h141E]=8'h29; mem['h141F]=8'hF1;
    mem['h1420]=8'hE3; mem['h1421]=8'h01; mem['h1422]=8'hCE; mem['h1423]=8'h13;
    mem['h1424]=8'hC5; mem['h1425]=8'h3D; mem['h1426]=8'hBE; mem['h1427]=8'h06;
    mem['h1428]=8'h00; mem['h1429]=8'hD0; mem['h142A]=8'h4F; mem['h142B]=8'h7E;
    mem['h142C]=8'h91; mem['h142D]=8'hBB; mem['h142E]=8'h47; mem['h142F]=8'hD8;
    mem['h1430]=8'h43; mem['h1431]=8'hC9; mem['h1432]=8'hCD; mem['h1433]=8'h9C;
    mem['h1434]=8'h13; mem['h1435]=8'hCA; mem['h1436]=8'h4F; mem['h1437]=8'h15;
    mem['h1438]=8'h5F; mem['h1439]=8'h23; mem['h143A]=8'h23; mem['h143B]=8'h7E;
    mem['h143C]=8'h23; mem['h143D]=8'h66; mem['h143E]=8'h6F; mem['h143F]=8'hE5;
    mem['h1440]=8'h19; mem['h1441]=8'h46; mem['h1442]=8'h72; mem['h1443]=8'hE3;
    mem['h1444]=8'hC5; mem['h1445]=8'h7E; mem['h1446]=8'hFE; mem['h1447]=8'h24;
    mem['h1448]=8'hC2; mem['h1449]=8'h50; mem['h144A]=8'h14; mem['h144B]=8'hCD;
    mem['h144C]=8'h7A; mem['h144D]=8'h1C; mem['h144E]=8'h18; mem['h144F]=8'h0D;
    mem['h1450]=8'hFE; mem['h1451]=8'h25; mem['h1452]=8'hC2; mem['h1453]=8'h5A;
    mem['h1454]=8'h14; mem['h1455]=8'hCD; mem['h1456]=8'hEA; mem['h1457]=8'h1C;
    mem['h1458]=8'h18; mem['h1459]=8'h03; mem['h145A]=8'hCD; mem['h145B]=8'h36;
    mem['h145C]=8'h18; mem['h145D]=8'hC1; mem['h145E]=8'hE1; mem['h145F]=8'h70;
    mem['h1460]=8'hC9; mem['h1461]=8'hEB; mem['h1462]=8'hCD; mem['h1463]=8'h56;
    mem['h1464]=8'h07; mem['h1465]=8'h29; mem['h1466]=8'hC1; mem['h1467]=8'hD1;
    mem['h1468]=8'hC5; mem['h1469]=8'h43; mem['h146A]=8'hC9; mem['h146B]=8'hCD;
    mem['h146C]=8'hB1; mem['h146D]=8'h14; mem['h146E]=8'h32; mem['h146F]=8'h84;
    mem['h1470]=8'h80; mem['h1471]=8'hCD; mem['h1472]=8'h83; mem['h1473]=8'h80;
    mem['h1474]=8'hC3; mem['h1475]=8'h17; mem['h1476]=8'h11; mem['h1477]=8'hCD;
    mem['h1478]=8'h9B; mem['h1479]=8'h14; mem['h147A]=8'hC3; mem['h147B]=8'h4B;
    mem['h147C]=8'h80; mem['h147D]=8'hCD; mem['h147E]=8'h9B; mem['h147F]=8'h14;
    mem['h1480]=8'hF5; mem['h1481]=8'h1E; mem['h1482]=8'h00; mem['h1483]=8'h2B;
    mem['h1484]=8'hCD; mem['h1485]=8'hE0; mem['h1486]=8'h08; mem['h1487]=8'hCA;
    mem['h1488]=8'h91; mem['h1489]=8'h14; mem['h148A]=8'hCD; mem['h148B]=8'h56;
    mem['h148C]=8'h07; mem['h148D]=8'h2C; mem['h148E]=8'hCD; mem['h148F]=8'hAE;
    mem['h1490]=8'h14; mem['h1491]=8'hC1; mem['h1492]=8'hCD; mem['h1493]=8'h83;
    mem['h1494]=8'h80; mem['h1495]=8'hAB; mem['h1496]=8'hA0; mem['h1497]=8'hCA;
    mem['h1498]=8'h92; mem['h1499]=8'h14; mem['h149A]=8'hC9; mem['h149B]=8'hCD;
    mem['h149C]=8'hAE; mem['h149D]=8'h14; mem['h149E]=8'h32; mem['h149F]=8'h84;
    mem['h14A0]=8'h80; mem['h14A1]=8'h32; mem['h14A2]=8'h4C; mem['h14A3]=8'h80;
    mem['h14A4]=8'hCD; mem['h14A5]=8'h56; mem['h14A6]=8'h07; mem['h14A7]=8'h2C;
    mem['h14A8]=8'hC3; mem['h14A9]=8'hAE; mem['h14AA]=8'h14; mem['h14AB]=8'hCD;
    mem['h14AC]=8'hE0; mem['h14AD]=8'h08; mem['h14AE]=8'hCD; mem['h14AF]=8'h4D;
    mem['h14B0]=8'h0D; mem['h14B1]=8'hCD; mem['h14B2]=8'h8C; mem['h14B3]=8'h09;
    mem['h14B4]=8'h7A; mem['h14B5]=8'hB7; mem['h14B6]=8'hC2; mem['h14B7]=8'hA7;
    mem['h14B8]=8'h09; mem['h14B9]=8'h2B; mem['h14BA]=8'hCD; mem['h14BB]=8'hE0;
    mem['h14BC]=8'h08; mem['h14BD]=8'h7B; mem['h14BE]=8'hC9; mem['h14BF]=8'hCD;
    mem['h14C0]=8'h92; mem['h14C1]=8'h09; mem['h14C2]=8'h1A; mem['h14C3]=8'hC3;
    mem['h14C4]=8'h17; mem['h14C5]=8'h11; mem['h14C6]=8'hCD; mem['h14C7]=8'h4D;
    mem['h14C8]=8'h0D; mem['h14C9]=8'hCD; mem['h14CA]=8'h92; mem['h14CB]=8'h09;
    mem['h14CC]=8'hD5; mem['h14CD]=8'hCD; mem['h14CE]=8'h56; mem['h14CF]=8'h07;
    mem['h14D0]=8'h2C; mem['h14D1]=8'hCD; mem['h14D2]=8'hAE; mem['h14D3]=8'h14;
    mem['h14D4]=8'hD1; mem['h14D5]=8'h12; mem['h14D6]=8'hC9; mem['h14D7]=8'h21;
    mem['h14D8]=8'hAD; mem['h14D9]=8'h19; mem['h14DA]=8'hCD; mem['h14DB]=8'h7E;
    mem['h14DC]=8'h17; mem['h14DD]=8'hC3; mem['h14DE]=8'hE9; mem['h14DF]=8'h14;
    mem['h14E0]=8'hCD; mem['h14E1]=8'h7E; mem['h14E2]=8'h17; mem['h14E3]=8'h21;
    mem['h14E4]=8'hC1; mem['h14E5]=8'hD1; mem['h14E6]=8'hCD; mem['h14E7]=8'h58;
    mem['h14E8]=8'h17; mem['h14E9]=8'h78; mem['h14EA]=8'hB7; mem['h14EB]=8'hC8;
    mem['h14EC]=8'h3A; mem['h14ED]=8'h2C; mem['h14EE]=8'h81; mem['h14EF]=8'hB7;
    mem['h14F0]=8'hCA; mem['h14F1]=8'h70; mem['h14F2]=8'h17; mem['h14F3]=8'h90;
    mem['h14F4]=8'hD2; mem['h14F5]=8'h03; mem['h14F6]=8'h15; mem['h14F7]=8'h2F;
    mem['h14F8]=8'h3C; mem['h14F9]=8'hEB; mem['h14FA]=8'hCD; mem['h14FB]=8'h60;
    mem['h14FC]=8'h17; mem['h14FD]=8'hEB; mem['h14FE]=8'hCD; mem['h14FF]=8'h70;
    mem['h1500]=8'h17; mem['h1501]=8'hC1; mem['h1502]=8'hD1; mem['h1503]=8'hFE;
    mem['h1504]=8'h19; mem['h1505]=8'hD0; mem['h1506]=8'hF5; mem['h1507]=8'hCD;
    mem['h1508]=8'h95; mem['h1509]=8'h17; mem['h150A]=8'h67; mem['h150B]=8'hF1;
    mem['h150C]=8'hCD; mem['h150D]=8'hAE; mem['h150E]=8'h15; mem['h150F]=8'hB4;
    mem['h1510]=8'h21; mem['h1511]=8'h29; mem['h1512]=8'h81; mem['h1513]=8'hF2;
    mem['h1514]=8'h29; mem['h1515]=8'h15; mem['h1516]=8'hCD; mem['h1517]=8'h8E;
    mem['h1518]=8'h15; mem['h1519]=8'hD2; mem['h151A]=8'h6F; mem['h151B]=8'h15;
    mem['h151C]=8'h23; mem['h151D]=8'h34; mem['h151E]=8'hCA; mem['h151F]=8'h97;
    mem['h1520]=8'h04; mem['h1521]=8'h2E; mem['h1522]=8'h01; mem['h1523]=8'hCD;
    mem['h1524]=8'hC4; mem['h1525]=8'h15; mem['h1526]=8'hC3; mem['h1527]=8'h6F;
    mem['h1528]=8'h15; mem['h1529]=8'hAF; mem['h152A]=8'h90; mem['h152B]=8'h47;
    mem['h152C]=8'h7E; mem['h152D]=8'h9B; mem['h152E]=8'h5F; mem['h152F]=8'h23;
    mem['h1530]=8'h7E; mem['h1531]=8'h9A; mem['h1532]=8'h57; mem['h1533]=8'h23;
    mem['h1534]=8'h7E; mem['h1535]=8'h99; mem['h1536]=8'h4F; mem['h1537]=8'hDC;
    mem['h1538]=8'h9A; mem['h1539]=8'h15; mem['h153A]=8'h68; mem['h153B]=8'h63;
    mem['h153C]=8'hAF; mem['h153D]=8'h47; mem['h153E]=8'h79; mem['h153F]=8'hB7;
    mem['h1540]=8'hC2; mem['h1541]=8'h5C; mem['h1542]=8'h15; mem['h1543]=8'h4A;
    mem['h1544]=8'h54; mem['h1545]=8'h65; mem['h1546]=8'h6F; mem['h1547]=8'h78;
    mem['h1548]=8'hD6; mem['h1549]=8'h08; mem['h154A]=8'hFE; mem['h154B]=8'hE0;
    mem['h154C]=8'hC2; mem['h154D]=8'h3D; mem['h154E]=8'h15; mem['h154F]=8'hAF;
    mem['h1550]=8'h32; mem['h1551]=8'h2C; mem['h1552]=8'h81; mem['h1553]=8'hC9;
    mem['h1554]=8'h05; mem['h1555]=8'h29; mem['h1556]=8'h7A; mem['h1557]=8'h17;
    mem['h1558]=8'h57; mem['h1559]=8'h79; mem['h155A]=8'h8F; mem['h155B]=8'h4F;
    mem['h155C]=8'hF2; mem['h155D]=8'h54; mem['h155E]=8'h15; mem['h155F]=8'h78;
    mem['h1560]=8'h5C; mem['h1561]=8'h45; mem['h1562]=8'hB7; mem['h1563]=8'hCA;
    mem['h1564]=8'h6F; mem['h1565]=8'h15; mem['h1566]=8'h21; mem['h1567]=8'h2C;
    mem['h1568]=8'h81; mem['h1569]=8'h86; mem['h156A]=8'h77; mem['h156B]=8'hD2;
    mem['h156C]=8'h4F; mem['h156D]=8'h15; mem['h156E]=8'hC8; mem['h156F]=8'h78;
    mem['h1570]=8'h21; mem['h1571]=8'h2C; mem['h1572]=8'h81; mem['h1573]=8'hB7;
    mem['h1574]=8'hFC; mem['h1575]=8'h81; mem['h1576]=8'h15; mem['h1577]=8'h46;
    mem['h1578]=8'h23; mem['h1579]=8'h7E; mem['h157A]=8'hE6; mem['h157B]=8'h80;
    mem['h157C]=8'hA9; mem['h157D]=8'h4F; mem['h157E]=8'hC3; mem['h157F]=8'h70;
    mem['h1580]=8'h17; mem['h1581]=8'h1C; mem['h1582]=8'hC0; mem['h1583]=8'h14;
    mem['h1584]=8'hC0; mem['h1585]=8'h0C; mem['h1586]=8'hC0; mem['h1587]=8'h0E;
    mem['h1588]=8'h80; mem['h1589]=8'h34; mem['h158A]=8'hC0; mem['h158B]=8'hC3;
    mem['h158C]=8'h97; mem['h158D]=8'h04; mem['h158E]=8'h7E; mem['h158F]=8'h83;
    mem['h1590]=8'h5F; mem['h1591]=8'h23; mem['h1592]=8'h7E; mem['h1593]=8'h8A;
    mem['h1594]=8'h57; mem['h1595]=8'h23; mem['h1596]=8'h7E; mem['h1597]=8'h89;
    mem['h1598]=8'h4F; mem['h1599]=8'hC9; mem['h159A]=8'h21; mem['h159B]=8'h2D;
    mem['h159C]=8'h81; mem['h159D]=8'h7E; mem['h159E]=8'h2F; mem['h159F]=8'h77;
    mem['h15A0]=8'hAF; mem['h15A1]=8'h6F; mem['h15A2]=8'h90; mem['h15A3]=8'h47;
    mem['h15A4]=8'h7D; mem['h15A5]=8'h9B; mem['h15A6]=8'h5F; mem['h15A7]=8'h7D;
    mem['h15A8]=8'h9A; mem['h15A9]=8'h57; mem['h15AA]=8'h7D; mem['h15AB]=8'h99;
    mem['h15AC]=8'h4F; mem['h15AD]=8'hC9; mem['h15AE]=8'h06; mem['h15AF]=8'h00;
    mem['h15B0]=8'hD6; mem['h15B1]=8'h08; mem['h15B2]=8'hDA; mem['h15B3]=8'hBD;
    mem['h15B4]=8'h15; mem['h15B5]=8'h43; mem['h15B6]=8'h5A; mem['h15B7]=8'h51;
    mem['h15B8]=8'h0E; mem['h15B9]=8'h00; mem['h15BA]=8'hC3; mem['h15BB]=8'hB0;
    mem['h15BC]=8'h15; mem['h15BD]=8'hC6; mem['h15BE]=8'h09; mem['h15BF]=8'h6F;
    mem['h15C0]=8'hAF; mem['h15C1]=8'h2D; mem['h15C2]=8'hC8; mem['h15C3]=8'h79;
    mem['h15C4]=8'h1F; mem['h15C5]=8'h4F; mem['h15C6]=8'h7A; mem['h15C7]=8'h1F;
    mem['h15C8]=8'h57; mem['h15C9]=8'h7B; mem['h15CA]=8'h1F; mem['h15CB]=8'h5F;
    mem['h15CC]=8'h78; mem['h15CD]=8'h1F; mem['h15CE]=8'h47; mem['h15CF]=8'hC3;
    mem['h15D0]=8'hC0; mem['h15D1]=8'h15; mem['h15D2]=8'h00; mem['h15D3]=8'h00;
    mem['h15D4]=8'h00; mem['h15D5]=8'h81; mem['h15D6]=8'h03; mem['h15D7]=8'hAA;
    mem['h15D8]=8'h56; mem['h15D9]=8'h19; mem['h15DA]=8'h80; mem['h15DB]=8'hF1;
    mem['h15DC]=8'h22; mem['h15DD]=8'h76; mem['h15DE]=8'h80; mem['h15DF]=8'h45;
    mem['h15E0]=8'hAA; mem['h15E1]=8'h38; mem['h15E2]=8'h82; mem['h15E3]=8'hCD;
    mem['h15E4]=8'h2F; mem['h15E5]=8'h17; mem['h15E6]=8'hB7; mem['h15E7]=8'hEA;
    mem['h15E8]=8'hA7; mem['h15E9]=8'h09; mem['h15EA]=8'h21; mem['h15EB]=8'h2C;
    mem['h15EC]=8'h81; mem['h15ED]=8'h7E; mem['h15EE]=8'h01; mem['h15EF]=8'h35;
    mem['h15F0]=8'h80; mem['h15F1]=8'h11; mem['h15F2]=8'hF3; mem['h15F3]=8'h04;
    mem['h15F4]=8'h90; mem['h15F5]=8'hF5; mem['h15F6]=8'h70; mem['h15F7]=8'hD5;
    mem['h15F8]=8'hC5; mem['h15F9]=8'hCD; mem['h15FA]=8'hE9; mem['h15FB]=8'h14;
    mem['h15FC]=8'hC1; mem['h15FD]=8'hD1; mem['h15FE]=8'h04; mem['h15FF]=8'hCD;
    mem['h1600]=8'h85; mem['h1601]=8'h16; mem['h1602]=8'h21; mem['h1603]=8'hD2;
    mem['h1604]=8'h15; mem['h1605]=8'hCD; mem['h1606]=8'hE0; mem['h1607]=8'h14;
    mem['h1608]=8'h21; mem['h1609]=8'hD6; mem['h160A]=8'h15; mem['h160B]=8'hCD;
    mem['h160C]=8'h77; mem['h160D]=8'h1A; mem['h160E]=8'h01; mem['h160F]=8'h80;
    mem['h1610]=8'h80; mem['h1611]=8'h11; mem['h1612]=8'h00; mem['h1613]=8'h00;
    mem['h1614]=8'hCD; mem['h1615]=8'hE9; mem['h1616]=8'h14; mem['h1617]=8'hF1;
    mem['h1618]=8'hCD; mem['h1619]=8'hAA; mem['h161A]=8'h18; mem['h161B]=8'h01;
    mem['h161C]=8'h31; mem['h161D]=8'h80; mem['h161E]=8'h11; mem['h161F]=8'h18;
    mem['h1620]=8'h72; mem['h1621]=8'h21; mem['h1622]=8'hC1; mem['h1623]=8'hD1;
    mem['h1624]=8'hCD; mem['h1625]=8'h2F; mem['h1626]=8'h17; mem['h1627]=8'hC8;
    mem['h1628]=8'h2E; mem['h1629]=8'h00; mem['h162A]=8'hCD; mem['h162B]=8'hED;
    mem['h162C]=8'h16; mem['h162D]=8'h79; mem['h162E]=8'h32; mem['h162F]=8'h3B;
    mem['h1630]=8'h81; mem['h1631]=8'hEB; mem['h1632]=8'h22; mem['h1633]=8'h3C;
    mem['h1634]=8'h81; mem['h1635]=8'h01; mem['h1636]=8'h00; mem['h1637]=8'h00;
    mem['h1638]=8'h50; mem['h1639]=8'h58; mem['h163A]=8'h21; mem['h163B]=8'h3A;
    mem['h163C]=8'h15; mem['h163D]=8'hE5; mem['h163E]=8'h21; mem['h163F]=8'h46;
    mem['h1640]=8'h16; mem['h1641]=8'hE5; mem['h1642]=8'hE5; mem['h1643]=8'h21;
    mem['h1644]=8'h29; mem['h1645]=8'h81; mem['h1646]=8'h7E; mem['h1647]=8'h23;
    mem['h1648]=8'hB7; mem['h1649]=8'hCA; mem['h164A]=8'h72; mem['h164B]=8'h16;
    mem['h164C]=8'hE5; mem['h164D]=8'h2E; mem['h164E]=8'h08; mem['h164F]=8'h1F;
    mem['h1650]=8'h67; mem['h1651]=8'h79; mem['h1652]=8'hD2; mem['h1653]=8'h60;
    mem['h1654]=8'h16; mem['h1655]=8'hE5; mem['h1656]=8'h2A; mem['h1657]=8'h3C;
    mem['h1658]=8'h81; mem['h1659]=8'h19; mem['h165A]=8'hEB; mem['h165B]=8'hE1;
    mem['h165C]=8'h3A; mem['h165D]=8'h3B; mem['h165E]=8'h81; mem['h165F]=8'h89;
    mem['h1660]=8'h1F; mem['h1661]=8'h4F; mem['h1662]=8'h7A; mem['h1663]=8'h1F;
    mem['h1664]=8'h57; mem['h1665]=8'h7B; mem['h1666]=8'h1F; mem['h1667]=8'h5F;
    mem['h1668]=8'h78; mem['h1669]=8'h1F; mem['h166A]=8'h47; mem['h166B]=8'h2D;
    mem['h166C]=8'h7C; mem['h166D]=8'hC2; mem['h166E]=8'h4F; mem['h166F]=8'h16;
    mem['h1670]=8'hE1; mem['h1671]=8'hC9; mem['h1672]=8'h43; mem['h1673]=8'h5A;
    mem['h1674]=8'h51; mem['h1675]=8'h4F; mem['h1676]=8'hC9; mem['h1677]=8'hCD;
    mem['h1678]=8'h60; mem['h1679]=8'h17; mem['h167A]=8'h01; mem['h167B]=8'h20;
    mem['h167C]=8'h84; mem['h167D]=8'h11; mem['h167E]=8'h00; mem['h167F]=8'h00;
    mem['h1680]=8'hCD; mem['h1681]=8'h70; mem['h1682]=8'h17; mem['h1683]=8'hC1;
    mem['h1684]=8'hD1; mem['h1685]=8'hCD; mem['h1686]=8'h2F; mem['h1687]=8'h17;
    mem['h1688]=8'hCA; mem['h1689]=8'h8B; mem['h168A]=8'h04; mem['h168B]=8'h2E;
    mem['h168C]=8'hFF; mem['h168D]=8'hCD; mem['h168E]=8'hED; mem['h168F]=8'h16;
    mem['h1690]=8'h34; mem['h1691]=8'h34; mem['h1692]=8'h2B; mem['h1693]=8'h7E;
    mem['h1694]=8'h32; mem['h1695]=8'h57; mem['h1696]=8'h80; mem['h1697]=8'h2B;
    mem['h1698]=8'h7E; mem['h1699]=8'h32; mem['h169A]=8'h53; mem['h169B]=8'h80;
    mem['h169C]=8'h2B; mem['h169D]=8'h7E; mem['h169E]=8'h32; mem['h169F]=8'h4F;
    mem['h16A0]=8'h80; mem['h16A1]=8'h41; mem['h16A2]=8'hEB; mem['h16A3]=8'hAF;
    mem['h16A4]=8'h4F; mem['h16A5]=8'h57; mem['h16A6]=8'h5F; mem['h16A7]=8'h32;
    mem['h16A8]=8'h5A; mem['h16A9]=8'h80; mem['h16AA]=8'hE5; mem['h16AB]=8'hC5;
    mem['h16AC]=8'h7D; mem['h16AD]=8'hCD; mem['h16AE]=8'h4E; mem['h16AF]=8'h80;
    mem['h16B0]=8'hDE; mem['h16B1]=8'h00; mem['h16B2]=8'h3F; mem['h16B3]=8'hD2;
    mem['h16B4]=8'hBD; mem['h16B5]=8'h16; mem['h16B6]=8'h32; mem['h16B7]=8'h5A;
    mem['h16B8]=8'h80; mem['h16B9]=8'hF1; mem['h16BA]=8'hF1; mem['h16BB]=8'h37;
    mem['h16BC]=8'hD2; mem['h16BD]=8'hC1; mem['h16BE]=8'hE1; mem['h16BF]=8'h79;
    mem['h16C0]=8'h3C; mem['h16C1]=8'h3D; mem['h16C2]=8'h1F; mem['h16C3]=8'hFA;
    mem['h16C4]=8'h70; mem['h16C5]=8'h15; mem['h16C6]=8'h17; mem['h16C7]=8'h7B;
    mem['h16C8]=8'h17; mem['h16C9]=8'h5F; mem['h16CA]=8'h7A; mem['h16CB]=8'h17;
    mem['h16CC]=8'h57; mem['h16CD]=8'h79; mem['h16CE]=8'h17; mem['h16CF]=8'h4F;
    mem['h16D0]=8'h29; mem['h16D1]=8'h78; mem['h16D2]=8'h17; mem['h16D3]=8'h47;
    mem['h16D4]=8'h3A; mem['h16D5]=8'h5A; mem['h16D6]=8'h80; mem['h16D7]=8'h17;
    mem['h16D8]=8'h32; mem['h16D9]=8'h5A; mem['h16DA]=8'h80; mem['h16DB]=8'h79;
    mem['h16DC]=8'hB2; mem['h16DD]=8'hB3; mem['h16DE]=8'hC2; mem['h16DF]=8'hAA;
    mem['h16E0]=8'h16; mem['h16E1]=8'hE5; mem['h16E2]=8'h21; mem['h16E3]=8'h2C;
    mem['h16E4]=8'h81; mem['h16E5]=8'h35; mem['h16E6]=8'hE1; mem['h16E7]=8'hC2;
    mem['h16E8]=8'hAA; mem['h16E9]=8'h16; mem['h16EA]=8'hC3; mem['h16EB]=8'h97;
    mem['h16EC]=8'h04; mem['h16ED]=8'h78; mem['h16EE]=8'hB7; mem['h16EF]=8'hCA;
    mem['h16F0]=8'h11; mem['h16F1]=8'h17; mem['h16F2]=8'h7D; mem['h16F3]=8'h21;
    mem['h16F4]=8'h2C; mem['h16F5]=8'h81; mem['h16F6]=8'hAE; mem['h16F7]=8'h80;
    mem['h16F8]=8'h47; mem['h16F9]=8'h1F; mem['h16FA]=8'hA8; mem['h16FB]=8'h78;
    mem['h16FC]=8'hF2; mem['h16FD]=8'h10; mem['h16FE]=8'h17; mem['h16FF]=8'hC6;
    mem['h1700]=8'h80; mem['h1701]=8'h77; mem['h1702]=8'hCA; mem['h1703]=8'h70;
    mem['h1704]=8'h16; mem['h1705]=8'hCD; mem['h1706]=8'h95; mem['h1707]=8'h17;
    mem['h1708]=8'h77; mem['h1709]=8'h2B; mem['h170A]=8'hC9; mem['h170B]=8'hCD;
    mem['h170C]=8'h2F; mem['h170D]=8'h17; mem['h170E]=8'h2F; mem['h170F]=8'hE1;
    mem['h1710]=8'hB7; mem['h1711]=8'hE1; mem['h1712]=8'hF2; mem['h1713]=8'h4F;
    mem['h1714]=8'h15; mem['h1715]=8'hC3; mem['h1716]=8'h97; mem['h1717]=8'h04;
    mem['h1718]=8'hCD; mem['h1719]=8'h7B; mem['h171A]=8'h17; mem['h171B]=8'h78;
    mem['h171C]=8'hB7; mem['h171D]=8'hC8; mem['h171E]=8'hC6; mem['h171F]=8'h02;
    mem['h1720]=8'hDA; mem['h1721]=8'h97; mem['h1722]=8'h04; mem['h1723]=8'h47;
    mem['h1724]=8'hCD; mem['h1725]=8'hE9; mem['h1726]=8'h14; mem['h1727]=8'h21;
    mem['h1728]=8'h2C; mem['h1729]=8'h81; mem['h172A]=8'h34; mem['h172B]=8'hC0;
    mem['h172C]=8'hC3; mem['h172D]=8'h97; mem['h172E]=8'h04; mem['h172F]=8'h3A;
    mem['h1730]=8'h2C; mem['h1731]=8'h81; mem['h1732]=8'hB7; mem['h1733]=8'hC8;
    mem['h1734]=8'h3A; mem['h1735]=8'h2B; mem['h1736]=8'h81; mem['h1737]=8'hFE;
    mem['h1738]=8'h2F; mem['h1739]=8'h17; mem['h173A]=8'h9F; mem['h173B]=8'hC0;
    mem['h173C]=8'h3C; mem['h173D]=8'hC9; mem['h173E]=8'hCD; mem['h173F]=8'h2F;
    mem['h1740]=8'h17; mem['h1741]=8'h06; mem['h1742]=8'h88; mem['h1743]=8'h11;
    mem['h1744]=8'h00; mem['h1745]=8'h00; mem['h1746]=8'h21; mem['h1747]=8'h2C;
    mem['h1748]=8'h81; mem['h1749]=8'h4F; mem['h174A]=8'h70; mem['h174B]=8'h06;
    mem['h174C]=8'h00; mem['h174D]=8'h23; mem['h174E]=8'h36; mem['h174F]=8'h80;
    mem['h1750]=8'h17; mem['h1751]=8'hC3; mem['h1752]=8'h37; mem['h1753]=8'h15;
    mem['h1754]=8'hCD; mem['h1755]=8'h2F; mem['h1756]=8'h17; mem['h1757]=8'hF0;
    mem['h1758]=8'h21; mem['h1759]=8'h2B; mem['h175A]=8'h81; mem['h175B]=8'h7E;
    mem['h175C]=8'hEE; mem['h175D]=8'h80; mem['h175E]=8'h77; mem['h175F]=8'hC9;
    mem['h1760]=8'hEB; mem['h1761]=8'h2A; mem['h1762]=8'h29; mem['h1763]=8'h81;
    mem['h1764]=8'hE3; mem['h1765]=8'hE5; mem['h1766]=8'h2A; mem['h1767]=8'h2B;
    mem['h1768]=8'h81; mem['h1769]=8'hE3; mem['h176A]=8'hE5; mem['h176B]=8'hEB;
    mem['h176C]=8'hC9; mem['h176D]=8'hCD; mem['h176E]=8'h7E; mem['h176F]=8'h17;
    mem['h1770]=8'hEB; mem['h1771]=8'h22; mem['h1772]=8'h29; mem['h1773]=8'h81;
    mem['h1774]=8'h60; mem['h1775]=8'h69; mem['h1776]=8'h22; mem['h1777]=8'h2B;
    mem['h1778]=8'h81; mem['h1779]=8'hEB; mem['h177A]=8'hC9; mem['h177B]=8'h21;
    mem['h177C]=8'h29; mem['h177D]=8'h81; mem['h177E]=8'h5E; mem['h177F]=8'h23;
    mem['h1780]=8'h56; mem['h1781]=8'h23; mem['h1782]=8'h4E; mem['h1783]=8'h23;
    mem['h1784]=8'h46; mem['h1785]=8'h23; mem['h1786]=8'hC9; mem['h1787]=8'h11;
    mem['h1788]=8'h29; mem['h1789]=8'h81; mem['h178A]=8'h06; mem['h178B]=8'h04;
    mem['h178C]=8'h1A; mem['h178D]=8'h77; mem['h178E]=8'h13; mem['h178F]=8'h23;
    mem['h1790]=8'h05; mem['h1791]=8'hC2; mem['h1792]=8'h8C; mem['h1793]=8'h17;
    mem['h1794]=8'hC9; mem['h1795]=8'h21; mem['h1796]=8'h2B; mem['h1797]=8'h81;
    mem['h1798]=8'h7E; mem['h1799]=8'h07; mem['h179A]=8'h37; mem['h179B]=8'h1F;
    mem['h179C]=8'h77; mem['h179D]=8'h3F; mem['h179E]=8'h1F; mem['h179F]=8'h23;
    mem['h17A0]=8'h23; mem['h17A1]=8'h77; mem['h17A2]=8'h79; mem['h17A3]=8'h07;
    mem['h17A4]=8'h37; mem['h17A5]=8'h1F; mem['h17A6]=8'h4F; mem['h17A7]=8'h1F;
    mem['h17A8]=8'hAE; mem['h17A9]=8'hC9; mem['h17AA]=8'h78; mem['h17AB]=8'hB7;
    mem['h17AC]=8'hCA; mem['h17AD]=8'h2F; mem['h17AE]=8'h17; mem['h17AF]=8'h21;
    mem['h17B0]=8'h38; mem['h17B1]=8'h17; mem['h17B2]=8'hE5; mem['h17B3]=8'hCD;
    mem['h17B4]=8'h2F; mem['h17B5]=8'h17; mem['h17B6]=8'h79; mem['h17B7]=8'hC8;
    mem['h17B8]=8'h21; mem['h17B9]=8'h2B; mem['h17BA]=8'h81; mem['h17BB]=8'hAE;
    mem['h17BC]=8'h79; mem['h17BD]=8'hF8; mem['h17BE]=8'hCD; mem['h17BF]=8'hC4;
    mem['h17C0]=8'h17; mem['h17C1]=8'h1F; mem['h17C2]=8'hA9; mem['h17C3]=8'hC9;
    mem['h17C4]=8'h23; mem['h17C5]=8'h78; mem['h17C6]=8'hBE; mem['h17C7]=8'hC0;
    mem['h17C8]=8'h2B; mem['h17C9]=8'h79; mem['h17CA]=8'hBE; mem['h17CB]=8'hC0;
    mem['h17CC]=8'h2B; mem['h17CD]=8'h7A; mem['h17CE]=8'hBE; mem['h17CF]=8'hC0;
    mem['h17D0]=8'h2B; mem['h17D1]=8'h7B; mem['h17D2]=8'h96; mem['h17D3]=8'hC0;
    mem['h17D4]=8'hE1; mem['h17D5]=8'hE1; mem['h17D6]=8'hC9; mem['h17D7]=8'h47;
    mem['h17D8]=8'h4F; mem['h17D9]=8'h57; mem['h17DA]=8'h5F; mem['h17DB]=8'hB7;
    mem['h17DC]=8'hC8; mem['h17DD]=8'hE5; mem['h17DE]=8'hCD; mem['h17DF]=8'h7B;
    mem['h17E0]=8'h17; mem['h17E1]=8'hCD; mem['h17E2]=8'h95; mem['h17E3]=8'h17;
    mem['h17E4]=8'hAE; mem['h17E5]=8'h67; mem['h17E6]=8'hFC; mem['h17E7]=8'hFB;
    mem['h17E8]=8'h17; mem['h17E9]=8'h3E; mem['h17EA]=8'h98; mem['h17EB]=8'h90;
    mem['h17EC]=8'hCD; mem['h17ED]=8'hAE; mem['h17EE]=8'h15; mem['h17EF]=8'h7C;
    mem['h17F0]=8'h17; mem['h17F1]=8'hDC; mem['h17F2]=8'h81; mem['h17F3]=8'h15;
    mem['h17F4]=8'h06; mem['h17F5]=8'h00; mem['h17F6]=8'hDC; mem['h17F7]=8'h9A;
    mem['h17F8]=8'h15; mem['h17F9]=8'hE1; mem['h17FA]=8'hC9; mem['h17FB]=8'h1B;
    mem['h17FC]=8'h7A; mem['h17FD]=8'hA3; mem['h17FE]=8'h3C; mem['h17FF]=8'hC0;
    mem['h1800]=8'h0B; mem['h1801]=8'hC9; mem['h1802]=8'h21; mem['h1803]=8'h2C;
    mem['h1804]=8'h81; mem['h1805]=8'h7E; mem['h1806]=8'hFE; mem['h1807]=8'h98;
    mem['h1808]=8'h3A; mem['h1809]=8'h29; mem['h180A]=8'h81; mem['h180B]=8'hD0;
    mem['h180C]=8'h7E; mem['h180D]=8'hCD; mem['h180E]=8'hD7; mem['h180F]=8'h17;
    mem['h1810]=8'h36; mem['h1811]=8'h98; mem['h1812]=8'h7B; mem['h1813]=8'hF5;
    mem['h1814]=8'h79; mem['h1815]=8'h17; mem['h1816]=8'hCD; mem['h1817]=8'h37;
    mem['h1818]=8'h15; mem['h1819]=8'hF1; mem['h181A]=8'hC9; mem['h181B]=8'h21;
    mem['h181C]=8'h00; mem['h181D]=8'h00; mem['h181E]=8'h78; mem['h181F]=8'hB1;
    mem['h1820]=8'hC8; mem['h1821]=8'h3E; mem['h1822]=8'h10; mem['h1823]=8'h29;
    mem['h1824]=8'hDA; mem['h1825]=8'h5B; mem['h1826]=8'h10; mem['h1827]=8'hEB;
    mem['h1828]=8'h29; mem['h1829]=8'hEB; mem['h182A]=8'hD2; mem['h182B]=8'h31;
    mem['h182C]=8'h18; mem['h182D]=8'h09; mem['h182E]=8'hDA; mem['h182F]=8'h5B;
    mem['h1830]=8'h10; mem['h1831]=8'h3D; mem['h1832]=8'hC2; mem['h1833]=8'h23;
    mem['h1834]=8'h18; mem['h1835]=8'hC9; mem['h1836]=8'hFE; mem['h1837]=8'h2D;
    mem['h1838]=8'hF5; mem['h1839]=8'hCA; mem['h183A]=8'h42; mem['h183B]=8'h18;
    mem['h183C]=8'hFE; mem['h183D]=8'h2B; mem['h183E]=8'hCA; mem['h183F]=8'h42;
    mem['h1840]=8'h18; mem['h1841]=8'h2B; mem['h1842]=8'hCD; mem['h1843]=8'h4F;
    mem['h1844]=8'h15; mem['h1845]=8'h47; mem['h1846]=8'h57; mem['h1847]=8'h5F;
    mem['h1848]=8'h2F; mem['h1849]=8'h4F; mem['h184A]=8'hCD; mem['h184B]=8'hE0;
    mem['h184C]=8'h08; mem['h184D]=8'hDA; mem['h184E]=8'h93; mem['h184F]=8'h18;
    mem['h1850]=8'hFE; mem['h1851]=8'h2E; mem['h1852]=8'hCA; mem['h1853]=8'h6E;
    mem['h1854]=8'h18; mem['h1855]=8'hFE; mem['h1856]=8'h45; mem['h1857]=8'hC2;
    mem['h1858]=8'h72; mem['h1859]=8'h18; mem['h185A]=8'hCD; mem['h185B]=8'hE0;
    mem['h185C]=8'h08; mem['h185D]=8'hCD; mem['h185E]=8'h86; mem['h185F]=8'h0E;
    mem['h1860]=8'hCD; mem['h1861]=8'hE0; mem['h1862]=8'h08; mem['h1863]=8'hDA;
    mem['h1864]=8'hB5; mem['h1865]=8'h18; mem['h1866]=8'h14; mem['h1867]=8'hC2;
    mem['h1868]=8'h72; mem['h1869]=8'h18; mem['h186A]=8'hAF; mem['h186B]=8'h93;
    mem['h186C]=8'h5F; mem['h186D]=8'h0C; mem['h186E]=8'h0C; mem['h186F]=8'hCA;
    mem['h1870]=8'h4A; mem['h1871]=8'h18; mem['h1872]=8'hE5; mem['h1873]=8'h7B;
    mem['h1874]=8'h90; mem['h1875]=8'hF4; mem['h1876]=8'h8B; mem['h1877]=8'h18;
    mem['h1878]=8'hF2; mem['h1879]=8'h81; mem['h187A]=8'h18; mem['h187B]=8'hF5;
    mem['h187C]=8'hCD; mem['h187D]=8'h77; mem['h187E]=8'h16; mem['h187F]=8'hF1;
    mem['h1880]=8'h3C; mem['h1881]=8'hC2; mem['h1882]=8'h75; mem['h1883]=8'h18;
    mem['h1884]=8'hD1; mem['h1885]=8'hF1; mem['h1886]=8'hCC; mem['h1887]=8'h58;
    mem['h1888]=8'h17; mem['h1889]=8'hEB; mem['h188A]=8'hC9; mem['h188B]=8'hC8;
    mem['h188C]=8'hF5; mem['h188D]=8'hCD; mem['h188E]=8'h18; mem['h188F]=8'h17;
    mem['h1890]=8'hF1; mem['h1891]=8'h3D; mem['h1892]=8'hC9; mem['h1893]=8'hD5;
    mem['h1894]=8'h57; mem['h1895]=8'h78; mem['h1896]=8'h89; mem['h1897]=8'h47;
    mem['h1898]=8'hC5; mem['h1899]=8'hE5; mem['h189A]=8'hD5; mem['h189B]=8'hCD;
    mem['h189C]=8'h18; mem['h189D]=8'h17; mem['h189E]=8'hF1; mem['h189F]=8'hD6;
    mem['h18A0]=8'h30; mem['h18A1]=8'hCD; mem['h18A2]=8'hAA; mem['h18A3]=8'h18;
    mem['h18A4]=8'hE1; mem['h18A5]=8'hC1; mem['h18A6]=8'hD1; mem['h18A7]=8'hC3;
    mem['h18A8]=8'h4A; mem['h18A9]=8'h18; mem['h18AA]=8'hCD; mem['h18AB]=8'h60;
    mem['h18AC]=8'h17; mem['h18AD]=8'hCD; mem['h18AE]=8'h41; mem['h18AF]=8'h17;
    mem['h18B0]=8'hC1; mem['h18B1]=8'hD1; mem['h18B2]=8'hC3; mem['h18B3]=8'hE9;
    mem['h18B4]=8'h14; mem['h18B5]=8'h7B; mem['h18B6]=8'h07; mem['h18B7]=8'h07;
    mem['h18B8]=8'h83; mem['h18B9]=8'h07; mem['h18BA]=8'h86; mem['h18BB]=8'hD6;
    mem['h18BC]=8'h30; mem['h18BD]=8'h5F; mem['h18BE]=8'hC3; mem['h18BF]=8'h60;
    mem['h18C0]=8'h18; mem['h18C1]=8'hE5; mem['h18C2]=8'h21; mem['h18C3]=8'h20;
    mem['h18C4]=8'h04; mem['h18C5]=8'hCD; mem['h18C6]=8'h26; mem['h18C7]=8'h12;
    mem['h18C8]=8'hE1; mem['h18C9]=8'hEB; mem['h18CA]=8'hAF; mem['h18CB]=8'h06;
    mem['h18CC]=8'h98; mem['h18CD]=8'hCD; mem['h18CE]=8'h46; mem['h18CF]=8'h17;
    mem['h18D0]=8'h21; mem['h18D1]=8'h25; mem['h18D2]=8'h12; mem['h18D3]=8'hE5;
    mem['h18D4]=8'h21; mem['h18D5]=8'h2E; mem['h18D6]=8'h81; mem['h18D7]=8'hE5;
    mem['h18D8]=8'hCD; mem['h18D9]=8'h2F; mem['h18DA]=8'h17; mem['h18DB]=8'h36;
    mem['h18DC]=8'h20; mem['h18DD]=8'hF2; mem['h18DE]=8'hE2; mem['h18DF]=8'h18;
    mem['h18E0]=8'h36; mem['h18E1]=8'h2D; mem['h18E2]=8'h23; mem['h18E3]=8'h36;
    mem['h18E4]=8'h30; mem['h18E5]=8'hCA; mem['h18E6]=8'h98; mem['h18E7]=8'h19;
    mem['h18E8]=8'hE5; mem['h18E9]=8'hFC; mem['h18EA]=8'h58; mem['h18EB]=8'h17;
    mem['h18EC]=8'hAF; mem['h18ED]=8'hF5; mem['h18EE]=8'hCD; mem['h18EF]=8'h9E;
    mem['h18F0]=8'h19; mem['h18F1]=8'h01; mem['h18F2]=8'h43; mem['h18F3]=8'h91;
    mem['h18F4]=8'h11; mem['h18F5]=8'hF8; mem['h18F6]=8'h4F; mem['h18F7]=8'hCD;
    mem['h18F8]=8'hAA; mem['h18F9]=8'h17; mem['h18FA]=8'hB7; mem['h18FB]=8'hE2;
    mem['h18FC]=8'h0F; mem['h18FD]=8'h19; mem['h18FE]=8'hF1; mem['h18FF]=8'hCD;
    mem['h1900]=8'h8C; mem['h1901]=8'h18; mem['h1902]=8'hF5; mem['h1903]=8'hC3;
    mem['h1904]=8'hF1; mem['h1905]=8'h18; mem['h1906]=8'hCD; mem['h1907]=8'h77;
    mem['h1908]=8'h16; mem['h1909]=8'hF1; mem['h190A]=8'h3C; mem['h190B]=8'hF5;
    mem['h190C]=8'hCD; mem['h190D]=8'h9E; mem['h190E]=8'h19; mem['h190F]=8'hCD;
    mem['h1910]=8'hD7; mem['h1911]=8'h14; mem['h1912]=8'h3C; mem['h1913]=8'hCD;
    mem['h1914]=8'hD7; mem['h1915]=8'h17; mem['h1916]=8'hCD; mem['h1917]=8'h70;
    mem['h1918]=8'h17; mem['h1919]=8'h01; mem['h191A]=8'h06; mem['h191B]=8'h03;
    mem['h191C]=8'hF1; mem['h191D]=8'h81; mem['h191E]=8'h3C; mem['h191F]=8'hFA;
    mem['h1920]=8'h2B; mem['h1921]=8'h19; mem['h1922]=8'hFE; mem['h1923]=8'h08;
    mem['h1924]=8'hD2; mem['h1925]=8'h2B; mem['h1926]=8'h19; mem['h1927]=8'h3C;
    mem['h1928]=8'h47; mem['h1929]=8'h3E; mem['h192A]=8'h02; mem['h192B]=8'h3D;
    mem['h192C]=8'h3D; mem['h192D]=8'hE1; mem['h192E]=8'hF5; mem['h192F]=8'h11;
    mem['h1930]=8'hB1; mem['h1931]=8'h19; mem['h1932]=8'h05; mem['h1933]=8'hC2;
    mem['h1934]=8'h3C; mem['h1935]=8'h19; mem['h1936]=8'h36; mem['h1937]=8'h2E;
    mem['h1938]=8'h23; mem['h1939]=8'h36; mem['h193A]=8'h30; mem['h193B]=8'h23;
    mem['h193C]=8'h05; mem['h193D]=8'h36; mem['h193E]=8'h2E; mem['h193F]=8'hCC;
    mem['h1940]=8'h85; mem['h1941]=8'h17; mem['h1942]=8'hC5; mem['h1943]=8'hE5;
    mem['h1944]=8'hD5; mem['h1945]=8'hCD; mem['h1946]=8'h7B; mem['h1947]=8'h17;
    mem['h1948]=8'hE1; mem['h1949]=8'h06; mem['h194A]=8'h2F; mem['h194B]=8'h04;
    mem['h194C]=8'h7B; mem['h194D]=8'h96; mem['h194E]=8'h5F; mem['h194F]=8'h23;
    mem['h1950]=8'h7A; mem['h1951]=8'h9E; mem['h1952]=8'h57; mem['h1953]=8'h23;
    mem['h1954]=8'h79; mem['h1955]=8'h9E; mem['h1956]=8'h4F; mem['h1957]=8'h2B;
    mem['h1958]=8'h2B; mem['h1959]=8'hD2; mem['h195A]=8'h4B; mem['h195B]=8'h19;
    mem['h195C]=8'hCD; mem['h195D]=8'h8E; mem['h195E]=8'h15; mem['h195F]=8'h23;
    mem['h1960]=8'hCD; mem['h1961]=8'h70; mem['h1962]=8'h17; mem['h1963]=8'hEB;
    mem['h1964]=8'hE1; mem['h1965]=8'h70; mem['h1966]=8'h23; mem['h1967]=8'hC1;
    mem['h1968]=8'h0D; mem['h1969]=8'hC2; mem['h196A]=8'h3C; mem['h196B]=8'h19;
    mem['h196C]=8'h05; mem['h196D]=8'hCA; mem['h196E]=8'h7C; mem['h196F]=8'h19;
    mem['h1970]=8'h2B; mem['h1971]=8'h7E; mem['h1972]=8'hFE; mem['h1973]=8'h30;
    mem['h1974]=8'hCA; mem['h1975]=8'h70; mem['h1976]=8'h19; mem['h1977]=8'hFE;
    mem['h1978]=8'h2E; mem['h1979]=8'hC4; mem['h197A]=8'h85; mem['h197B]=8'h17;
    mem['h197C]=8'hF1; mem['h197D]=8'hCA; mem['h197E]=8'h9B; mem['h197F]=8'h19;
    mem['h1980]=8'h36; mem['h1981]=8'h45; mem['h1982]=8'h23; mem['h1983]=8'h36;
    mem['h1984]=8'h2B; mem['h1985]=8'hF2; mem['h1986]=8'h8C; mem['h1987]=8'h19;
    mem['h1988]=8'h36; mem['h1989]=8'h2D; mem['h198A]=8'h2F; mem['h198B]=8'h3C;
    mem['h198C]=8'h06; mem['h198D]=8'h2F; mem['h198E]=8'h04; mem['h198F]=8'hD6;
    mem['h1990]=8'h0A; mem['h1991]=8'hD2; mem['h1992]=8'h8E; mem['h1993]=8'h19;
    mem['h1994]=8'hC6; mem['h1995]=8'h3A; mem['h1996]=8'h23; mem['h1997]=8'h70;
    mem['h1998]=8'h23; mem['h1999]=8'h77; mem['h199A]=8'h23; mem['h199B]=8'h71;
    mem['h199C]=8'hE1; mem['h199D]=8'hC9; mem['h199E]=8'h01; mem['h199F]=8'h74;
    mem['h19A0]=8'h94; mem['h19A1]=8'h11; mem['h19A2]=8'hF7; mem['h19A3]=8'h23;
    mem['h19A4]=8'hCD; mem['h19A5]=8'hAA; mem['h19A6]=8'h17; mem['h19A7]=8'hB7;
    mem['h19A8]=8'hE1; mem['h19A9]=8'hE2; mem['h19AA]=8'h06; mem['h19AB]=8'h19;
    mem['h19AC]=8'hE9; mem['h19AD]=8'h00; mem['h19AE]=8'h00; mem['h19AF]=8'h00;
    mem['h19B0]=8'h80; mem['h19B1]=8'hA0; mem['h19B2]=8'h86; mem['h19B3]=8'h01;
    mem['h19B4]=8'h10; mem['h19B5]=8'h27; mem['h19B6]=8'h00; mem['h19B7]=8'hE8;
    mem['h19B8]=8'h03; mem['h19B9]=8'h00; mem['h19BA]=8'h64; mem['h19BB]=8'h00;
    mem['h19BC]=8'h00; mem['h19BD]=8'h0A; mem['h19BE]=8'h00; mem['h19BF]=8'h00;
    mem['h19C0]=8'h01; mem['h19C1]=8'h00; mem['h19C2]=8'h00; mem['h19C3]=8'h21;
    mem['h19C4]=8'h58; mem['h19C5]=8'h17; mem['h19C6]=8'hE3; mem['h19C7]=8'hE9;
    mem['h19C8]=8'hCD; mem['h19C9]=8'h60; mem['h19CA]=8'h17; mem['h19CB]=8'h21;
    mem['h19CC]=8'hAD; mem['h19CD]=8'h19; mem['h19CE]=8'hCD; mem['h19CF]=8'h6D;
    mem['h19D0]=8'h17; mem['h19D1]=8'hC1; mem['h19D2]=8'hD1; mem['h19D3]=8'hCD;
    mem['h19D4]=8'h2F; mem['h19D5]=8'h17; mem['h19D6]=8'h78; mem['h19D7]=8'hCA;
    mem['h19D8]=8'h16; mem['h19D9]=8'h1A; mem['h19DA]=8'hF2; mem['h19DB]=8'hE1;
    mem['h19DC]=8'h19; mem['h19DD]=8'hB7; mem['h19DE]=8'hCA; mem['h19DF]=8'h8B;
    mem['h19E0]=8'h04; mem['h19E1]=8'hB7; mem['h19E2]=8'hCA; mem['h19E3]=8'h50;
    mem['h19E4]=8'h15; mem['h19E5]=8'hD5; mem['h19E6]=8'hC5; mem['h19E7]=8'h79;
    mem['h19E8]=8'hF6; mem['h19E9]=8'h7F; mem['h19EA]=8'hCD; mem['h19EB]=8'h7B;
    mem['h19EC]=8'h17; mem['h19ED]=8'hF2; mem['h19EE]=8'hFE; mem['h19EF]=8'h19;
    mem['h19F0]=8'hD5; mem['h19F1]=8'hC5; mem['h19F2]=8'hCD; mem['h19F3]=8'h02;
    mem['h19F4]=8'h18; mem['h19F5]=8'hC1; mem['h19F6]=8'hD1; mem['h19F7]=8'hF5;
    mem['h19F8]=8'hCD; mem['h19F9]=8'hAA; mem['h19FA]=8'h17; mem['h19FB]=8'hE1;
    mem['h19FC]=8'h7C; mem['h19FD]=8'h1F; mem['h19FE]=8'hE1; mem['h19FF]=8'h22;
    mem['h1A00]=8'h2B; mem['h1A01]=8'h81; mem['h1A02]=8'hE1; mem['h1A03]=8'h22;
    mem['h1A04]=8'h29; mem['h1A05]=8'h81; mem['h1A06]=8'hDC; mem['h1A07]=8'hC3;
    mem['h1A08]=8'h19; mem['h1A09]=8'hCC; mem['h1A0A]=8'h58; mem['h1A0B]=8'h17;
    mem['h1A0C]=8'hD5; mem['h1A0D]=8'hC5; mem['h1A0E]=8'hCD; mem['h1A0F]=8'hE3;
    mem['h1A10]=8'h15; mem['h1A11]=8'hC1; mem['h1A12]=8'hD1; mem['h1A13]=8'hCD;
    mem['h1A14]=8'h24; mem['h1A15]=8'h16; mem['h1A16]=8'hCD; mem['h1A17]=8'h60;
    mem['h1A18]=8'h17; mem['h1A19]=8'h01; mem['h1A1A]=8'h38; mem['h1A1B]=8'h81;
    mem['h1A1C]=8'h11; mem['h1A1D]=8'h3B; mem['h1A1E]=8'hAA; mem['h1A1F]=8'hCD;
    mem['h1A20]=8'h24; mem['h1A21]=8'h16; mem['h1A22]=8'h3A; mem['h1A23]=8'h2C;
    mem['h1A24]=8'h81; mem['h1A25]=8'hFE; mem['h1A26]=8'h88; mem['h1A27]=8'hD2;
    mem['h1A28]=8'h0B; mem['h1A29]=8'h17; mem['h1A2A]=8'hCD; mem['h1A2B]=8'h02;
    mem['h1A2C]=8'h18; mem['h1A2D]=8'hC6; mem['h1A2E]=8'h80; mem['h1A2F]=8'hC6;
    mem['h1A30]=8'h02; mem['h1A31]=8'hDA; mem['h1A32]=8'h0B; mem['h1A33]=8'h17;
    mem['h1A34]=8'hF5; mem['h1A35]=8'h21; mem['h1A36]=8'hD2; mem['h1A37]=8'h15;
    mem['h1A38]=8'hCD; mem['h1A39]=8'hDA; mem['h1A3A]=8'h14; mem['h1A3B]=8'hCD;
    mem['h1A3C]=8'h1B; mem['h1A3D]=8'h16; mem['h1A3E]=8'hF1; mem['h1A3F]=8'hC1;
    mem['h1A40]=8'hD1; mem['h1A41]=8'hF5; mem['h1A42]=8'hCD; mem['h1A43]=8'hE6;
    mem['h1A44]=8'h14; mem['h1A45]=8'hCD; mem['h1A46]=8'h58; mem['h1A47]=8'h17;
    mem['h1A48]=8'h21; mem['h1A49]=8'h56; mem['h1A4A]=8'h1A; mem['h1A4B]=8'hCD;
    mem['h1A4C]=8'h86; mem['h1A4D]=8'h1A; mem['h1A4E]=8'h11; mem['h1A4F]=8'h00;
    mem['h1A50]=8'h00; mem['h1A51]=8'hC1; mem['h1A52]=8'h4A; mem['h1A53]=8'hC3;
    mem['h1A54]=8'h24; mem['h1A55]=8'h16; mem['h1A56]=8'h08; mem['h1A57]=8'h40;
    mem['h1A58]=8'h2E; mem['h1A59]=8'h94; mem['h1A5A]=8'h74; mem['h1A5B]=8'h70;
    mem['h1A5C]=8'h4F; mem['h1A5D]=8'h2E; mem['h1A5E]=8'h77; mem['h1A5F]=8'h6E;
    mem['h1A60]=8'h02; mem['h1A61]=8'h88; mem['h1A62]=8'h7A; mem['h1A63]=8'hE6;
    mem['h1A64]=8'hA0; mem['h1A65]=8'h2A; mem['h1A66]=8'h7C; mem['h1A67]=8'h50;
    mem['h1A68]=8'hAA; mem['h1A69]=8'hAA; mem['h1A6A]=8'h7E; mem['h1A6B]=8'hFF;
    mem['h1A6C]=8'hFF; mem['h1A6D]=8'h7F; mem['h1A6E]=8'h7F; mem['h1A6F]=8'h00;
    mem['h1A70]=8'h00; mem['h1A71]=8'h80; mem['h1A72]=8'h81; mem['h1A73]=8'h00;
    mem['h1A74]=8'h00; mem['h1A75]=8'h00; mem['h1A76]=8'h81; mem['h1A77]=8'hCD;
    mem['h1A78]=8'h60; mem['h1A79]=8'h17; mem['h1A7A]=8'h11; mem['h1A7B]=8'h22;
    mem['h1A7C]=8'h16; mem['h1A7D]=8'hD5; mem['h1A7E]=8'hE5; mem['h1A7F]=8'hCD;
    mem['h1A80]=8'h7B; mem['h1A81]=8'h17; mem['h1A82]=8'hCD; mem['h1A83]=8'h24;
    mem['h1A84]=8'h16; mem['h1A85]=8'hE1; mem['h1A86]=8'hCD; mem['h1A87]=8'h60;
    mem['h1A88]=8'h17; mem['h1A89]=8'h7E; mem['h1A8A]=8'h23; mem['h1A8B]=8'hCD;
    mem['h1A8C]=8'h6D; mem['h1A8D]=8'h17; mem['h1A8E]=8'h06; mem['h1A8F]=8'hF1;
    mem['h1A90]=8'hC1; mem['h1A91]=8'hD1; mem['h1A92]=8'h3D; mem['h1A93]=8'hC8;
    mem['h1A94]=8'hD5; mem['h1A95]=8'hC5; mem['h1A96]=8'hF5; mem['h1A97]=8'hE5;
    mem['h1A98]=8'hCD; mem['h1A99]=8'h24; mem['h1A9A]=8'h16; mem['h1A9B]=8'hE1;
    mem['h1A9C]=8'hCD; mem['h1A9D]=8'h7E; mem['h1A9E]=8'h17; mem['h1A9F]=8'hE5;
    mem['h1AA0]=8'hCD; mem['h1AA1]=8'hE9; mem['h1AA2]=8'h14; mem['h1AA3]=8'hE1;
    mem['h1AA4]=8'hC3; mem['h1AA5]=8'h8F; mem['h1AA6]=8'h1A; mem['h1AA7]=8'hCD;
    mem['h1AA8]=8'h2F; mem['h1AA9]=8'h17; mem['h1AAA]=8'h21; mem['h1AAB]=8'h5E;
    mem['h1AAC]=8'h80; mem['h1AAD]=8'hFA; mem['h1AAE]=8'h08; mem['h1AAF]=8'h1B;
    mem['h1AB0]=8'h21; mem['h1AB1]=8'h7F; mem['h1AB2]=8'h80; mem['h1AB3]=8'hCD;
    mem['h1AB4]=8'h6D; mem['h1AB5]=8'h17; mem['h1AB6]=8'h21; mem['h1AB7]=8'h5E;
    mem['h1AB8]=8'h80; mem['h1AB9]=8'hC8; mem['h1ABA]=8'h86; mem['h1ABB]=8'hE6;
    mem['h1ABC]=8'h07; mem['h1ABD]=8'h06; mem['h1ABE]=8'h00; mem['h1ABF]=8'h77;
    mem['h1AC0]=8'h23; mem['h1AC1]=8'h87; mem['h1AC2]=8'h87; mem['h1AC3]=8'h4F;
    mem['h1AC4]=8'h09; mem['h1AC5]=8'hCD; mem['h1AC6]=8'h7E; mem['h1AC7]=8'h17;
    mem['h1AC8]=8'hCD; mem['h1AC9]=8'h24; mem['h1ACA]=8'h16; mem['h1ACB]=8'h3A;
    mem['h1ACC]=8'h5D; mem['h1ACD]=8'h80; mem['h1ACE]=8'h3C; mem['h1ACF]=8'hE6;
    mem['h1AD0]=8'h03; mem['h1AD1]=8'h06; mem['h1AD2]=8'h00; mem['h1AD3]=8'hFE;
    mem['h1AD4]=8'h01; mem['h1AD5]=8'h88; mem['h1AD6]=8'h32; mem['h1AD7]=8'h5D;
    mem['h1AD8]=8'h80; mem['h1AD9]=8'h21; mem['h1ADA]=8'h0C; mem['h1ADB]=8'h1B;
    mem['h1ADC]=8'h87; mem['h1ADD]=8'h87; mem['h1ADE]=8'h4F; mem['h1ADF]=8'h09;
    mem['h1AE0]=8'hCD; mem['h1AE1]=8'hDA; mem['h1AE2]=8'h14; mem['h1AE3]=8'hCD;
    mem['h1AE4]=8'h7B; mem['h1AE5]=8'h17; mem['h1AE6]=8'h7B; mem['h1AE7]=8'h59;
    mem['h1AE8]=8'hEE; mem['h1AE9]=8'h4F; mem['h1AEA]=8'h4F; mem['h1AEB]=8'h36;
    mem['h1AEC]=8'h80; mem['h1AED]=8'h2B; mem['h1AEE]=8'h46; mem['h1AEF]=8'h36;
    mem['h1AF0]=8'h80; mem['h1AF1]=8'h21; mem['h1AF2]=8'h5C; mem['h1AF3]=8'h80;
    mem['h1AF4]=8'h34; mem['h1AF5]=8'h7E; mem['h1AF6]=8'hD6; mem['h1AF7]=8'hAB;
    mem['h1AF8]=8'hC2; mem['h1AF9]=8'hFF; mem['h1AFA]=8'h1A; mem['h1AFB]=8'h77;
    mem['h1AFC]=8'h0C; mem['h1AFD]=8'h15; mem['h1AFE]=8'h1C; mem['h1AFF]=8'hCD;
    mem['h1B00]=8'h3A; mem['h1B01]=8'h15; mem['h1B02]=8'h21; mem['h1B03]=8'h7F;
    mem['h1B04]=8'h80; mem['h1B05]=8'hC3; mem['h1B06]=8'h87; mem['h1B07]=8'h17;
    mem['h1B08]=8'h77; mem['h1B09]=8'h2B; mem['h1B0A]=8'h77; mem['h1B0B]=8'h2B;
    mem['h1B0C]=8'h77; mem['h1B0D]=8'hC3; mem['h1B0E]=8'hE3; mem['h1B0F]=8'h1A;
    mem['h1B10]=8'h68; mem['h1B11]=8'hB1; mem['h1B12]=8'h46; mem['h1B13]=8'h68;
    mem['h1B14]=8'h99; mem['h1B15]=8'hE9; mem['h1B16]=8'h92; mem['h1B17]=8'h69;
    mem['h1B18]=8'h10; mem['h1B19]=8'hD1; mem['h1B1A]=8'h75; mem['h1B1B]=8'h68;
    mem['h1B1C]=8'h21; mem['h1B1D]=8'h66; mem['h1B1E]=8'h1B; mem['h1B1F]=8'hCD;
    mem['h1B20]=8'hDA; mem['h1B21]=8'h14; mem['h1B22]=8'hCD; mem['h1B23]=8'h60;
    mem['h1B24]=8'h17; mem['h1B25]=8'h01; mem['h1B26]=8'h49; mem['h1B27]=8'h83;
    mem['h1B28]=8'h11; mem['h1B29]=8'hDB; mem['h1B2A]=8'h0F; mem['h1B2B]=8'hCD;
    mem['h1B2C]=8'h70; mem['h1B2D]=8'h17; mem['h1B2E]=8'hC1; mem['h1B2F]=8'hD1;
    mem['h1B30]=8'hCD; mem['h1B31]=8'h85; mem['h1B32]=8'h16; mem['h1B33]=8'hCD;
    mem['h1B34]=8'h60; mem['h1B35]=8'h17; mem['h1B36]=8'hCD; mem['h1B37]=8'h02;
    mem['h1B38]=8'h18; mem['h1B39]=8'hC1; mem['h1B3A]=8'hD1; mem['h1B3B]=8'hCD;
    mem['h1B3C]=8'hE6; mem['h1B3D]=8'h14; mem['h1B3E]=8'h21; mem['h1B3F]=8'h6A;
    mem['h1B40]=8'h1B; mem['h1B41]=8'hCD; mem['h1B42]=8'hE0; mem['h1B43]=8'h14;
    mem['h1B44]=8'hCD; mem['h1B45]=8'h2F; mem['h1B46]=8'h17; mem['h1B47]=8'h37;
    mem['h1B48]=8'hF2; mem['h1B49]=8'h52; mem['h1B4A]=8'h1B; mem['h1B4B]=8'hCD;
    mem['h1B4C]=8'hD7; mem['h1B4D]=8'h14; mem['h1B4E]=8'hCD; mem['h1B4F]=8'h2F;
    mem['h1B50]=8'h17; mem['h1B51]=8'hB7; mem['h1B52]=8'hF5; mem['h1B53]=8'hF4;
    mem['h1B54]=8'h58; mem['h1B55]=8'h17; mem['h1B56]=8'h21; mem['h1B57]=8'h6A;
    mem['h1B58]=8'h1B; mem['h1B59]=8'hCD; mem['h1B5A]=8'hDA; mem['h1B5B]=8'h14;
    mem['h1B5C]=8'hF1; mem['h1B5D]=8'hD4; mem['h1B5E]=8'h58; mem['h1B5F]=8'h17;
    mem['h1B60]=8'h21; mem['h1B61]=8'h6E; mem['h1B62]=8'h1B; mem['h1B63]=8'hC3;
    mem['h1B64]=8'h77; mem['h1B65]=8'h1A; mem['h1B66]=8'hDB; mem['h1B67]=8'h0F;
    mem['h1B68]=8'h49; mem['h1B69]=8'h81; mem['h1B6A]=8'h00; mem['h1B6B]=8'h00;
    mem['h1B6C]=8'h00; mem['h1B6D]=8'h7F; mem['h1B6E]=8'h05; mem['h1B6F]=8'hBA;
    mem['h1B70]=8'hD7; mem['h1B71]=8'h1E; mem['h1B72]=8'h86; mem['h1B73]=8'h64;
    mem['h1B74]=8'h26; mem['h1B75]=8'h99; mem['h1B76]=8'h87; mem['h1B77]=8'h58;
    mem['h1B78]=8'h34; mem['h1B79]=8'h23; mem['h1B7A]=8'h87; mem['h1B7B]=8'hE0;
    mem['h1B7C]=8'h5D; mem['h1B7D]=8'hA5; mem['h1B7E]=8'h86; mem['h1B7F]=8'hDA;
    mem['h1B80]=8'h0F; mem['h1B81]=8'h49; mem['h1B82]=8'h83; mem['h1B83]=8'hCD;
    mem['h1B84]=8'h60; mem['h1B85]=8'h17; mem['h1B86]=8'hCD; mem['h1B87]=8'h22;
    mem['h1B88]=8'h1B; mem['h1B89]=8'hC1; mem['h1B8A]=8'hE1; mem['h1B8B]=8'hCD;
    mem['h1B8C]=8'h60; mem['h1B8D]=8'h17; mem['h1B8E]=8'hEB; mem['h1B8F]=8'hCD;
    mem['h1B90]=8'h70; mem['h1B91]=8'h17; mem['h1B92]=8'hCD; mem['h1B93]=8'h1C;
    mem['h1B94]=8'h1B; mem['h1B95]=8'hC3; mem['h1B96]=8'h83; mem['h1B97]=8'h16;
    mem['h1B98]=8'hCD; mem['h1B99]=8'h2F; mem['h1B9A]=8'h17; mem['h1B9B]=8'hFC;
    mem['h1B9C]=8'hC3; mem['h1B9D]=8'h19; mem['h1B9E]=8'hFC; mem['h1B9F]=8'h58;
    mem['h1BA0]=8'h17; mem['h1BA1]=8'h3A; mem['h1BA2]=8'h2C; mem['h1BA3]=8'h81;
    mem['h1BA4]=8'hFE; mem['h1BA5]=8'h81; mem['h1BA6]=8'hDA; mem['h1BA7]=8'hB5;
    mem['h1BA8]=8'h1B; mem['h1BA9]=8'h01; mem['h1BAA]=8'h00; mem['h1BAB]=8'h81;
    mem['h1BAC]=8'h51; mem['h1BAD]=8'h59; mem['h1BAE]=8'hCD; mem['h1BAF]=8'h85;
    mem['h1BB0]=8'h16; mem['h1BB1]=8'h21; mem['h1BB2]=8'hE0; mem['h1BB3]=8'h14;
    mem['h1BB4]=8'hE5; mem['h1BB5]=8'h21; mem['h1BB6]=8'hBF; mem['h1BB7]=8'h1B;
    mem['h1BB8]=8'hCD; mem['h1BB9]=8'h77; mem['h1BBA]=8'h1A; mem['h1BBB]=8'h21;
    mem['h1BBC]=8'h66; mem['h1BBD]=8'h1B; mem['h1BBE]=8'hC9; mem['h1BBF]=8'h09;
    mem['h1BC0]=8'h4A; mem['h1BC1]=8'hD7; mem['h1BC2]=8'h3B; mem['h1BC3]=8'h78;
    mem['h1BC4]=8'h02; mem['h1BC5]=8'h6E; mem['h1BC6]=8'h84; mem['h1BC7]=8'h7B;
    mem['h1BC8]=8'hFE; mem['h1BC9]=8'hC1; mem['h1BCA]=8'h2F; mem['h1BCB]=8'h7C;
    mem['h1BCC]=8'h74; mem['h1BCD]=8'h31; mem['h1BCE]=8'h9A; mem['h1BCF]=8'h7D;
    mem['h1BD0]=8'h84; mem['h1BD1]=8'h3D; mem['h1BD2]=8'h5A; mem['h1BD3]=8'h7D;
    mem['h1BD4]=8'hC8; mem['h1BD5]=8'h7F; mem['h1BD6]=8'h91; mem['h1BD7]=8'h7E;
    mem['h1BD8]=8'hE4; mem['h1BD9]=8'hBB; mem['h1BDA]=8'h4C; mem['h1BDB]=8'h7E;
    mem['h1BDC]=8'h6C; mem['h1BDD]=8'hAA; mem['h1BDE]=8'hAA; mem['h1BDF]=8'h7F;
    mem['h1BE0]=8'h00; mem['h1BE1]=8'h00; mem['h1BE2]=8'h00; mem['h1BE3]=8'h81;
    mem['h1BE4]=8'hC9; mem['h1BE5]=8'hD7; mem['h1BE6]=8'hC9; mem['h1BE7]=8'h3E;
    mem['h1BE8]=8'h0C; mem['h1BE9]=8'hC3; mem['h1BEA]=8'h1D; mem['h1BEB]=8'h1D;
    mem['h1BEC]=8'hCD; mem['h1BED]=8'hAE; mem['h1BEE]=8'h14; mem['h1BEF]=8'h7B;
    mem['h1BF0]=8'h32; mem['h1BF1]=8'h87; mem['h1BF2]=8'h80; mem['h1BF3]=8'hC9;
    mem['h1BF4]=8'hCD; mem['h1BF5]=8'h4D; mem['h1BF6]=8'h0D; mem['h1BF7]=8'hCD;
    mem['h1BF8]=8'h92; mem['h1BF9]=8'h09; mem['h1BFA]=8'hED; mem['h1BFB]=8'h53;
    mem['h1BFC]=8'h8B; mem['h1BFD]=8'h80; mem['h1BFE]=8'hED; mem['h1BFF]=8'h53;
    mem['h1C00]=8'h8D; mem['h1C01]=8'h80; mem['h1C02]=8'hC9; mem['h1C03]=8'hCD;
    mem['h1C04]=8'h92; mem['h1C05]=8'h09; mem['h1C06]=8'hD5; mem['h1C07]=8'hE1;
    mem['h1C08]=8'h46; mem['h1C09]=8'h23; mem['h1C0A]=8'h7E; mem['h1C0B]=8'hC3;
    mem['h1C0C]=8'h08; mem['h1C0D]=8'h11; mem['h1C0E]=8'hCD; mem['h1C0F]=8'h4D;
    mem['h1C10]=8'h0D; mem['h1C11]=8'hCD; mem['h1C12]=8'h92; mem['h1C13]=8'h09;
    mem['h1C14]=8'hD5; mem['h1C15]=8'hCD; mem['h1C16]=8'h56; mem['h1C17]=8'h07;
    mem['h1C18]=8'h2C; mem['h1C19]=8'hCD; mem['h1C1A]=8'h4D; mem['h1C1B]=8'h0D;
    mem['h1C1C]=8'hCD; mem['h1C1D]=8'h92; mem['h1C1E]=8'h09; mem['h1C1F]=8'hE3;
    mem['h1C20]=8'h73; mem['h1C21]=8'h23; mem['h1C22]=8'h72; mem['h1C23]=8'hE1;
    mem['h1C24]=8'hC9; mem['h1C25]=8'hCD; mem['h1C26]=8'h50; mem['h1C27]=8'h0D;
    mem['h1C28]=8'hCD; mem['h1C29]=8'h92; mem['h1C2A]=8'h09; mem['h1C2B]=8'hC5;
    mem['h1C2C]=8'h21; mem['h1C2D]=8'h2E; mem['h1C2E]=8'h81; mem['h1C2F]=8'h7A;
    mem['h1C30]=8'hFE; mem['h1C31]=8'h00; mem['h1C32]=8'h28; mem['h1C33]=8'h0C;
    mem['h1C34]=8'hCD; mem['h1C35]=8'h5D; mem['h1C36]=8'h1C; mem['h1C37]=8'h78;
    mem['h1C38]=8'hFE; mem['h1C39]=8'h30; mem['h1C3A]=8'h28; mem['h1C3B]=8'h02;
    mem['h1C3C]=8'h70; mem['h1C3D]=8'h23; mem['h1C3E]=8'h71; mem['h1C3F]=8'h23;
    mem['h1C40]=8'h7B; mem['h1C41]=8'hCD; mem['h1C42]=8'h5D; mem['h1C43]=8'h1C;
    mem['h1C44]=8'h7A; mem['h1C45]=8'hFE; mem['h1C46]=8'h00; mem['h1C47]=8'h20;
    mem['h1C48]=8'h05; mem['h1C49]=8'h78; mem['h1C4A]=8'hFE; mem['h1C4B]=8'h30;
    mem['h1C4C]=8'h28; mem['h1C4D]=8'h02; mem['h1C4E]=8'h70; mem['h1C4F]=8'h23;
    mem['h1C50]=8'h71; mem['h1C51]=8'h23; mem['h1C52]=8'hAF; mem['h1C53]=8'h77;
    mem['h1C54]=8'h23; mem['h1C55]=8'h77; mem['h1C56]=8'hC1; mem['h1C57]=8'h21;
    mem['h1C58]=8'h2E; mem['h1C59]=8'h81; mem['h1C5A]=8'hC3; mem['h1C5B]=8'hB6;
    mem['h1C5C]=8'h11; mem['h1C5D]=8'h47; mem['h1C5E]=8'hE6; mem['h1C5F]=8'h0F;
    mem['h1C60]=8'hFE; mem['h1C61]=8'h0A; mem['h1C62]=8'h38; mem['h1C63]=8'h02;
    mem['h1C64]=8'hC6; mem['h1C65]=8'h07; mem['h1C66]=8'hC6; mem['h1C67]=8'h30;
    mem['h1C68]=8'h4F; mem['h1C69]=8'h78; mem['h1C6A]=8'h0F; mem['h1C6B]=8'h0F;
    mem['h1C6C]=8'h0F; mem['h1C6D]=8'h0F; mem['h1C6E]=8'hE6; mem['h1C6F]=8'h0F;
    mem['h1C70]=8'hFE; mem['h1C71]=8'h0A; mem['h1C72]=8'h38; mem['h1C73]=8'h02;
    mem['h1C74]=8'hC6; mem['h1C75]=8'h07; mem['h1C76]=8'hC6; mem['h1C77]=8'h30;
    mem['h1C78]=8'h47; mem['h1C79]=8'hC9; mem['h1C7A]=8'hEB; mem['h1C7B]=8'h21;
    mem['h1C7C]=8'h00; mem['h1C7D]=8'h00; mem['h1C7E]=8'hCD; mem['h1C7F]=8'h93;
    mem['h1C80]=8'h1C; mem['h1C81]=8'hDA; mem['h1C82]=8'hB3; mem['h1C83]=8'h1C;
    mem['h1C84]=8'h18; mem['h1C85]=8'h05; mem['h1C86]=8'hCD; mem['h1C87]=8'h93;
    mem['h1C88]=8'h1C; mem['h1C89]=8'h38; mem['h1C8A]=8'h1F; mem['h1C8B]=8'h29;
    mem['h1C8C]=8'h29; mem['h1C8D]=8'h29; mem['h1C8E]=8'h29; mem['h1C8F]=8'hB5;
    mem['h1C90]=8'h6F; mem['h1C91]=8'h18; mem['h1C92]=8'hF3; mem['h1C93]=8'h13;
    mem['h1C94]=8'h1A; mem['h1C95]=8'hFE; mem['h1C96]=8'h20; mem['h1C97]=8'hCA;
    mem['h1C98]=8'h93; mem['h1C99]=8'h1C; mem['h1C9A]=8'hD6; mem['h1C9B]=8'h30;
    mem['h1C9C]=8'hD8; mem['h1C9D]=8'hFE; mem['h1C9E]=8'h0A; mem['h1C9F]=8'h38;
    mem['h1CA0]=8'h05; mem['h1CA1]=8'hD6; mem['h1CA2]=8'h07; mem['h1CA3]=8'hFE;
    mem['h1CA4]=8'h0A; mem['h1CA5]=8'hD8; mem['h1CA6]=8'hFE; mem['h1CA7]=8'h10;
    mem['h1CA8]=8'h3F; mem['h1CA9]=8'hC9; mem['h1CAA]=8'hEB; mem['h1CAB]=8'h7A;
    mem['h1CAC]=8'h4B; mem['h1CAD]=8'hE5; mem['h1CAE]=8'hCD; mem['h1CAF]=8'h07;
    mem['h1CB0]=8'h11; mem['h1CB1]=8'hE1; mem['h1CB2]=8'hC9; mem['h1CB3]=8'h1E;
    mem['h1CB4]=8'h26; mem['h1CB5]=8'hC3; mem['h1CB6]=8'h9C; mem['h1CB7]=8'h04;
    mem['h1CB8]=8'hCD; mem['h1CB9]=8'h50; mem['h1CBA]=8'h0D; mem['h1CBB]=8'hCD;
    mem['h1CBC]=8'h92; mem['h1CBD]=8'h09; mem['h1CBE]=8'hC5; mem['h1CBF]=8'h21;
    mem['h1CC0]=8'h2E; mem['h1CC1]=8'h81; mem['h1CC2]=8'h06; mem['h1CC3]=8'h11;
    mem['h1CC4]=8'h05; mem['h1CC5]=8'h78; mem['h1CC6]=8'hFE; mem['h1CC7]=8'h01;
    mem['h1CC8]=8'h28; mem['h1CC9]=8'h08; mem['h1CCA]=8'hCB; mem['h1CCB]=8'h13;
    mem['h1CCC]=8'hCB; mem['h1CCD]=8'h12; mem['h1CCE]=8'h30; mem['h1CCF]=8'hF4;
    mem['h1CD0]=8'h18; mem['h1CD1]=8'h04; mem['h1CD2]=8'hCB; mem['h1CD3]=8'h13;
    mem['h1CD4]=8'hCB; mem['h1CD5]=8'h12; mem['h1CD6]=8'h3E; mem['h1CD7]=8'h30;
    mem['h1CD8]=8'hCE; mem['h1CD9]=8'h00; mem['h1CDA]=8'h77; mem['h1CDB]=8'h23;
    mem['h1CDC]=8'h05; mem['h1CDD]=8'h20; mem['h1CDE]=8'hF3; mem['h1CDF]=8'hAF;
    mem['h1CE0]=8'h77; mem['h1CE1]=8'h23; mem['h1CE2]=8'h77; mem['h1CE3]=8'hC1;
    mem['h1CE4]=8'h21; mem['h1CE5]=8'h2E; mem['h1CE6]=8'h81; mem['h1CE7]=8'hC3;
    mem['h1CE8]=8'hB6; mem['h1CE9]=8'h11; mem['h1CEA]=8'hEB; mem['h1CEB]=8'h21;
    mem['h1CEC]=8'h00; mem['h1CED]=8'h00; mem['h1CEE]=8'hCD; mem['h1CEF]=8'h07;
    mem['h1CF0]=8'h1D; mem['h1CF1]=8'hDA; mem['h1CF2]=8'h15; mem['h1CF3]=8'h1D;
    mem['h1CF4]=8'hD6; mem['h1CF5]=8'h30; mem['h1CF6]=8'h29; mem['h1CF7]=8'hB5;
    mem['h1CF8]=8'h6F; mem['h1CF9]=8'hCD; mem['h1CFA]=8'h07; mem['h1CFB]=8'h1D;
    mem['h1CFC]=8'h30; mem['h1CFD]=8'hF6; mem['h1CFE]=8'hEB; mem['h1CFF]=8'h7A;
    mem['h1D00]=8'h4B; mem['h1D01]=8'hE5; mem['h1D02]=8'hCD; mem['h1D03]=8'h07;
    mem['h1D04]=8'h11; mem['h1D05]=8'hE1; mem['h1D06]=8'hC9; mem['h1D07]=8'h13;
    mem['h1D08]=8'h1A; mem['h1D09]=8'hFE; mem['h1D0A]=8'h20; mem['h1D0B]=8'hCA;
    mem['h1D0C]=8'h07; mem['h1D0D]=8'h1D; mem['h1D0E]=8'hFE; mem['h1D0F]=8'h30;
    mem['h1D10]=8'hD8; mem['h1D11]=8'hFE; mem['h1D12]=8'h32; mem['h1D13]=8'h3F;
    mem['h1D14]=8'hC9; mem['h1D15]=8'h1E; mem['h1D16]=8'h28; mem['h1D17]=8'hC3;
    mem['h1D18]=8'h9C; mem['h1D19]=8'h04; mem['h1D1A]=8'hC3; mem['h1D1B]=8'hE1;
    mem['h1D1C]=8'h00; mem['h1D1D]=8'hC3; mem['h1D1E]=8'h08; mem['h1D1F]=8'h00;
    mem['h1D20]=8'hC3; mem['h1D21]=8'h00; mem['h1D22]=8'h00; mem['h1D23]=8'h3E;
    mem['h1D24]=8'h00; mem['h1D25]=8'h32; mem['h1D26]=8'h92; mem['h1D27]=8'h80;
    mem['h1D28]=8'hC3; mem['h1D29]=8'hE8; mem['h1D2A]=8'h00; mem['h1D2B]=8'hF5;
    mem['h1D2C]=8'hA0; mem['h1D2D]=8'hC1; mem['h1D2E]=8'hB8; mem['h1D2F]=8'h3E;
    mem['h1D30]=8'h00; mem['h1D31]=8'hC9; mem['h1D32]=8'hCD; mem['h1D33]=8'h61;
    mem['h1D34]=8'h07; mem['h1D35]=8'hC3; mem['h1D36]=8'h88; mem['h1D37]=8'h0B;
    mem['h1D38]=8'hFF; mem['h1D39]=8'hFF; mem['h1D3A]=8'hFF; mem['h1D3B]=8'hFF;
    mem['h1D3C]=8'hFF; mem['h1D3D]=8'hFF; mem['h1D3E]=8'hFF; mem['h1D3F]=8'hFF;
    mem['h1D40]=8'hFF; mem['h1D41]=8'hFF; mem['h1D42]=8'hFF; mem['h1D43]=8'hFF;
    mem['h1D44]=8'hFF; mem['h1D45]=8'hFF; mem['h1D46]=8'hFF; mem['h1D47]=8'hFF;
    mem['h1D48]=8'hFF; mem['h1D49]=8'hFF; mem['h1D4A]=8'hFF; mem['h1D4B]=8'hFF;
    mem['h1D4C]=8'hFF; mem['h1D4D]=8'hFF; mem['h1D4E]=8'hFF; mem['h1D4F]=8'hFF;
    mem['h1D50]=8'hFF; mem['h1D51]=8'hFF; mem['h1D52]=8'hFF; mem['h1D53]=8'hFF;
    mem['h1D54]=8'hFF; mem['h1D55]=8'hFF; mem['h1D56]=8'hFF; mem['h1D57]=8'hFF;
    mem['h1D58]=8'hFF; mem['h1D59]=8'hFF; mem['h1D5A]=8'hFF; mem['h1D5B]=8'hFF;
    mem['h1D5C]=8'hFF; mem['h1D5D]=8'hFF; mem['h1D5E]=8'hFF; mem['h1D5F]=8'hFF;
    mem['h1D60]=8'hFF; mem['h1D61]=8'hFF; mem['h1D62]=8'hFF; mem['h1D63]=8'hFF;
    mem['h1D64]=8'hFF; mem['h1D65]=8'hFF; mem['h1D66]=8'hFF; mem['h1D67]=8'hFF;
    mem['h1D68]=8'hFF; mem['h1D69]=8'hFF; mem['h1D6A]=8'hFF; mem['h1D6B]=8'hFF;
    mem['h1D6C]=8'hFF; mem['h1D6D]=8'hFF; mem['h1D6E]=8'hFF; mem['h1D6F]=8'hFF;
    mem['h1D70]=8'hFF; mem['h1D71]=8'hFF; mem['h1D72]=8'hFF; mem['h1D73]=8'hFF;
    mem['h1D74]=8'hFF; mem['h1D75]=8'hFF; mem['h1D76]=8'hFF; mem['h1D77]=8'hFF;
    mem['h1D78]=8'hFF; mem['h1D79]=8'hFF; mem['h1D7A]=8'hFF; mem['h1D7B]=8'hFF;
    mem['h1D7C]=8'hFF; mem['h1D7D]=8'hFF; mem['h1D7E]=8'hFF; mem['h1D7F]=8'hFF;
    mem['h1D80]=8'hFF; mem['h1D81]=8'hFF; mem['h1D82]=8'hFF; mem['h1D83]=8'hFF;
    mem['h1D84]=8'hFF; mem['h1D85]=8'hFF; mem['h1D86]=8'hFF; mem['h1D87]=8'hFF;
    mem['h1D88]=8'hFF; mem['h1D89]=8'hFF; mem['h1D8A]=8'hFF; mem['h1D8B]=8'hFF;
    mem['h1D8C]=8'hFF; mem['h1D8D]=8'hFF; mem['h1D8E]=8'hFF; mem['h1D8F]=8'hFF;
    mem['h1D90]=8'hFF; mem['h1D91]=8'hFF; mem['h1D92]=8'hFF; mem['h1D93]=8'hFF;
    mem['h1D94]=8'hFF; mem['h1D95]=8'hFF; mem['h1D96]=8'hFF; mem['h1D97]=8'hFF;
    mem['h1D98]=8'hFF; mem['h1D99]=8'hFF; mem['h1D9A]=8'hFF; mem['h1D9B]=8'hFF;
    mem['h1D9C]=8'hFF; mem['h1D9D]=8'hFF; mem['h1D9E]=8'hFF; mem['h1D9F]=8'hFF;
    mem['h1DA0]=8'hFF; mem['h1DA1]=8'hFF; mem['h1DA2]=8'hFF; mem['h1DA3]=8'hFF;
    mem['h1DA4]=8'hFF; mem['h1DA5]=8'hFF; mem['h1DA6]=8'hFF; mem['h1DA7]=8'hFF;
    mem['h1DA8]=8'hFF; mem['h1DA9]=8'hFF; mem['h1DAA]=8'hFF; mem['h1DAB]=8'hFF;
    mem['h1DAC]=8'hFF; mem['h1DAD]=8'hFF; mem['h1DAE]=8'hFF; mem['h1DAF]=8'hFF;
    mem['h1DB0]=8'hFF; mem['h1DB1]=8'hFF; mem['h1DB2]=8'hFF; mem['h1DB3]=8'hFF;
    mem['h1DB4]=8'hFF; mem['h1DB5]=8'hFF; mem['h1DB6]=8'hFF; mem['h1DB7]=8'hFF;
    mem['h1DB8]=8'hFF; mem['h1DB9]=8'hFF; mem['h1DBA]=8'hFF; mem['h1DBB]=8'hFF;
    mem['h1DBC]=8'hFF; mem['h1DBD]=8'hFF; mem['h1DBE]=8'hFF; mem['h1DBF]=8'hFF;
    mem['h1DC0]=8'hFF; mem['h1DC1]=8'hFF; mem['h1DC2]=8'hFF; mem['h1DC3]=8'hFF;
    mem['h1DC4]=8'hFF; mem['h1DC5]=8'hFF; mem['h1DC6]=8'hFF; mem['h1DC7]=8'hFF;
    mem['h1DC8]=8'hFF; mem['h1DC9]=8'hFF; mem['h1DCA]=8'hFF; mem['h1DCB]=8'hFF;
    mem['h1DCC]=8'hFF; mem['h1DCD]=8'hFF; mem['h1DCE]=8'hFF; mem['h1DCF]=8'hFF;
    mem['h1DD0]=8'hFF; mem['h1DD1]=8'hFF; mem['h1DD2]=8'hFF; mem['h1DD3]=8'hFF;
    mem['h1DD4]=8'hFF; mem['h1DD5]=8'hFF; mem['h1DD6]=8'hFF; mem['h1DD7]=8'hFF;
    mem['h1DD8]=8'hFF; mem['h1DD9]=8'hFF; mem['h1DDA]=8'hFF; mem['h1DDB]=8'hFF;
    mem['h1DDC]=8'hFF; mem['h1DDD]=8'hFF; mem['h1DDE]=8'hFF; mem['h1DDF]=8'hFF;
    mem['h1DE0]=8'hFF; mem['h1DE1]=8'hFF; mem['h1DE2]=8'hFF; mem['h1DE3]=8'hFF;
    mem['h1DE4]=8'hFF; mem['h1DE5]=8'hFF; mem['h1DE6]=8'hFF; mem['h1DE7]=8'hFF;
    mem['h1DE8]=8'hFF; mem['h1DE9]=8'hFF; mem['h1DEA]=8'hFF; mem['h1DEB]=8'hFF;
    mem['h1DEC]=8'hFF; mem['h1DED]=8'hFF; mem['h1DEE]=8'hFF; mem['h1DEF]=8'hFF;
    mem['h1DF0]=8'hFF; mem['h1DF1]=8'hFF; mem['h1DF2]=8'hFF; mem['h1DF3]=8'hFF;
    mem['h1DF4]=8'hFF; mem['h1DF5]=8'hFF; mem['h1DF6]=8'hFF; mem['h1DF7]=8'hFF;
    mem['h1DF8]=8'hFF; mem['h1DF9]=8'hFF; mem['h1DFA]=8'hFF; mem['h1DFB]=8'hFF;
    mem['h1DFC]=8'hFF; mem['h1DFD]=8'hFF; mem['h1DFE]=8'hFF; mem['h1DFF]=8'hFF;
    mem['h1E00]=8'hFF; mem['h1E01]=8'hFF; mem['h1E02]=8'hFF; mem['h1E03]=8'hFF;
    mem['h1E04]=8'hFF; mem['h1E05]=8'hFF; mem['h1E06]=8'hFF; mem['h1E07]=8'hFF;
    mem['h1E08]=8'hFF; mem['h1E09]=8'hFF; mem['h1E0A]=8'hFF; mem['h1E0B]=8'hFF;
    mem['h1E0C]=8'hFF; mem['h1E0D]=8'hFF; mem['h1E0E]=8'hFF; mem['h1E0F]=8'hFF;
    mem['h1E10]=8'hFF; mem['h1E11]=8'hFF; mem['h1E12]=8'hFF; mem['h1E13]=8'hFF;
    mem['h1E14]=8'hFF; mem['h1E15]=8'hFF; mem['h1E16]=8'hFF; mem['h1E17]=8'hFF;
    mem['h1E18]=8'hFF; mem['h1E19]=8'hFF; mem['h1E1A]=8'hFF; mem['h1E1B]=8'hFF;
    mem['h1E1C]=8'hFF; mem['h1E1D]=8'hFF; mem['h1E1E]=8'hFF; mem['h1E1F]=8'hFF;
    mem['h1E20]=8'hFF; mem['h1E21]=8'hFF; mem['h1E22]=8'hFF; mem['h1E23]=8'hFF;
    mem['h1E24]=8'hFF; mem['h1E25]=8'hFF; mem['h1E26]=8'hFF; mem['h1E27]=8'hFF;
    mem['h1E28]=8'hFF; mem['h1E29]=8'hFF; mem['h1E2A]=8'hFF; mem['h1E2B]=8'hFF;
    mem['h1E2C]=8'hFF; mem['h1E2D]=8'hFF; mem['h1E2E]=8'hFF; mem['h1E2F]=8'hFF;
    mem['h1E30]=8'hFF; mem['h1E31]=8'hFF; mem['h1E32]=8'hFF; mem['h1E33]=8'hFF;
    mem['h1E34]=8'hFF; mem['h1E35]=8'hFF; mem['h1E36]=8'hFF; mem['h1E37]=8'hFF;
    mem['h1E38]=8'hFF; mem['h1E39]=8'hFF; mem['h1E3A]=8'hFF; mem['h1E3B]=8'hFF;
    mem['h1E3C]=8'hFF; mem['h1E3D]=8'hFF; mem['h1E3E]=8'hFF; mem['h1E3F]=8'hFF;
    mem['h1E40]=8'hFF; mem['h1E41]=8'hFF; mem['h1E42]=8'hFF; mem['h1E43]=8'hFF;
    mem['h1E44]=8'hFF; mem['h1E45]=8'hFF; mem['h1E46]=8'hFF; mem['h1E47]=8'hFF;
    mem['h1E48]=8'hFF; mem['h1E49]=8'hFF; mem['h1E4A]=8'hFF; mem['h1E4B]=8'hFF;
    mem['h1E4C]=8'hFF; mem['h1E4D]=8'hFF; mem['h1E4E]=8'hFF; mem['h1E4F]=8'hFF;
    mem['h1E50]=8'hFF; mem['h1E51]=8'hFF; mem['h1E52]=8'hFF; mem['h1E53]=8'hFF;
    mem['h1E54]=8'hFF; mem['h1E55]=8'hFF; mem['h1E56]=8'hFF; mem['h1E57]=8'hFF;
    mem['h1E58]=8'hFF; mem['h1E59]=8'hFF; mem['h1E5A]=8'hFF; mem['h1E5B]=8'hFF;
    mem['h1E5C]=8'hFF; mem['h1E5D]=8'hFF; mem['h1E5E]=8'hFF; mem['h1E5F]=8'hFF;
    mem['h1E60]=8'hFF; mem['h1E61]=8'hFF; mem['h1E62]=8'hFF; mem['h1E63]=8'hFF;
    mem['h1E64]=8'hFF; mem['h1E65]=8'hFF; mem['h1E66]=8'hFF; mem['h1E67]=8'hFF;
    mem['h1E68]=8'hFF; mem['h1E69]=8'hFF; mem['h1E6A]=8'hFF; mem['h1E6B]=8'hFF;
    mem['h1E6C]=8'hFF; mem['h1E6D]=8'hFF; mem['h1E6E]=8'hFF; mem['h1E6F]=8'hFF;
    mem['h1E70]=8'hFF; mem['h1E71]=8'hFF; mem['h1E72]=8'hFF; mem['h1E73]=8'hFF;
    mem['h1E74]=8'hFF; mem['h1E75]=8'hFF; mem['h1E76]=8'hFF; mem['h1E77]=8'hFF;
    mem['h1E78]=8'hFF; mem['h1E79]=8'hFF; mem['h1E7A]=8'hFF; mem['h1E7B]=8'hFF;
    mem['h1E7C]=8'hFF; mem['h1E7D]=8'hFF; mem['h1E7E]=8'hFF; mem['h1E7F]=8'hFF;
    mem['h1E80]=8'hFF; mem['h1E81]=8'hFF; mem['h1E82]=8'hFF; mem['h1E83]=8'hFF;
    mem['h1E84]=8'hFF; mem['h1E85]=8'hFF; mem['h1E86]=8'hFF; mem['h1E87]=8'hFF;
    mem['h1E88]=8'hFF; mem['h1E89]=8'hFF; mem['h1E8A]=8'hFF; mem['h1E8B]=8'hFF;
    mem['h1E8C]=8'hFF; mem['h1E8D]=8'hFF; mem['h1E8E]=8'hFF; mem['h1E8F]=8'hFF;
    mem['h1E90]=8'hFF; mem['h1E91]=8'hFF; mem['h1E92]=8'hFF; mem['h1E93]=8'hFF;
    mem['h1E94]=8'hFF; mem['h1E95]=8'hFF; mem['h1E96]=8'hFF; mem['h1E97]=8'hFF;
    mem['h1E98]=8'hFF; mem['h1E99]=8'hFF; mem['h1E9A]=8'hFF; mem['h1E9B]=8'hFF;
    mem['h1E9C]=8'hFF; mem['h1E9D]=8'hFF; mem['h1E9E]=8'hFF; mem['h1E9F]=8'hFF;
    mem['h1EA0]=8'hFF; mem['h1EA1]=8'hFF; mem['h1EA2]=8'hFF; mem['h1EA3]=8'hFF;
    mem['h1EA4]=8'hFF; mem['h1EA5]=8'hFF; mem['h1EA6]=8'hFF; mem['h1EA7]=8'hFF;
    mem['h1EA8]=8'hFF; mem['h1EA9]=8'hFF; mem['h1EAA]=8'hFF; mem['h1EAB]=8'hFF;
    mem['h1EAC]=8'hFF; mem['h1EAD]=8'hFF; mem['h1EAE]=8'hFF; mem['h1EAF]=8'hFF;
    mem['h1EB0]=8'hFF; mem['h1EB1]=8'hFF; mem['h1EB2]=8'hFF; mem['h1EB3]=8'hFF;
    mem['h1EB4]=8'hFF; mem['h1EB5]=8'hFF; mem['h1EB6]=8'hFF; mem['h1EB7]=8'hFF;
    mem['h1EB8]=8'hFF; mem['h1EB9]=8'hFF; mem['h1EBA]=8'hFF; mem['h1EBB]=8'hFF;
    mem['h1EBC]=8'hFF; mem['h1EBD]=8'hFF; mem['h1EBE]=8'hFF; mem['h1EBF]=8'hFF;
    mem['h1EC0]=8'hFF; mem['h1EC1]=8'hFF; mem['h1EC2]=8'hFF; mem['h1EC3]=8'hFF;
    mem['h1EC4]=8'hFF; mem['h1EC5]=8'hFF; mem['h1EC6]=8'hFF; mem['h1EC7]=8'hFF;
    mem['h1EC8]=8'hFF; mem['h1EC9]=8'hFF; mem['h1ECA]=8'hFF; mem['h1ECB]=8'hFF;
    mem['h1ECC]=8'hFF; mem['h1ECD]=8'hFF; mem['h1ECE]=8'hFF; mem['h1ECF]=8'hFF;
    mem['h1ED0]=8'hFF; mem['h1ED1]=8'hFF; mem['h1ED2]=8'hFF; mem['h1ED3]=8'hFF;
    mem['h1ED4]=8'hFF; mem['h1ED5]=8'hFF; mem['h1ED6]=8'hFF; mem['h1ED7]=8'hFF;
    mem['h1ED8]=8'hFF; mem['h1ED9]=8'hFF; mem['h1EDA]=8'hFF; mem['h1EDB]=8'hFF;
    mem['h1EDC]=8'hFF; mem['h1EDD]=8'hFF; mem['h1EDE]=8'hFF; mem['h1EDF]=8'hFF;
    mem['h1EE0]=8'hFF; mem['h1EE1]=8'hFF; mem['h1EE2]=8'hFF; mem['h1EE3]=8'hFF;
    mem['h1EE4]=8'hFF; mem['h1EE5]=8'hFF; mem['h1EE6]=8'hFF; mem['h1EE7]=8'hFF;
    mem['h1EE8]=8'hFF; mem['h1EE9]=8'hFF; mem['h1EEA]=8'hFF; mem['h1EEB]=8'hFF;
    mem['h1EEC]=8'hFF; mem['h1EED]=8'hFF; mem['h1EEE]=8'hFF; mem['h1EEF]=8'hFF;
    mem['h1EF0]=8'hFF; mem['h1EF1]=8'hFF; mem['h1EF2]=8'hFF; mem['h1EF3]=8'hFF;
    mem['h1EF4]=8'hFF; mem['h1EF5]=8'hFF; mem['h1EF6]=8'hFF; mem['h1EF7]=8'hFF;
    mem['h1EF8]=8'hFF; mem['h1EF9]=8'hFF; mem['h1EFA]=8'hFF; mem['h1EFB]=8'hFF;
    mem['h1EFC]=8'hFF; mem['h1EFD]=8'hFF; mem['h1EFE]=8'hFF; mem['h1EFF]=8'hFF;
    mem['h1F00]=8'hFF; mem['h1F01]=8'hFF; mem['h1F02]=8'hFF; mem['h1F03]=8'hFF;
    mem['h1F04]=8'hFF; mem['h1F05]=8'hFF; mem['h1F06]=8'hFF; mem['h1F07]=8'hFF;
    mem['h1F08]=8'hFF; mem['h1F09]=8'hFF; mem['h1F0A]=8'hFF; mem['h1F0B]=8'hFF;
    mem['h1F0C]=8'hFF; mem['h1F0D]=8'hFF; mem['h1F0E]=8'hFF; mem['h1F0F]=8'hFF;
    mem['h1F10]=8'hFF; mem['h1F11]=8'hFF; mem['h1F12]=8'hFF; mem['h1F13]=8'hFF;
    mem['h1F14]=8'hFF; mem['h1F15]=8'hFF; mem['h1F16]=8'hFF; mem['h1F17]=8'hFF;
    mem['h1F18]=8'hFF; mem['h1F19]=8'hFF; mem['h1F1A]=8'hFF; mem['h1F1B]=8'hFF;
    mem['h1F1C]=8'hFF; mem['h1F1D]=8'hFF; mem['h1F1E]=8'hFF; mem['h1F1F]=8'hFF;
    mem['h1F20]=8'hFF; mem['h1F21]=8'hFF; mem['h1F22]=8'hFF; mem['h1F23]=8'hFF;
    mem['h1F24]=8'hFF; mem['h1F25]=8'hFF; mem['h1F26]=8'hFF; mem['h1F27]=8'hFF;
    mem['h1F28]=8'hFF; mem['h1F29]=8'hFF; mem['h1F2A]=8'hFF; mem['h1F2B]=8'hFF;
    mem['h1F2C]=8'hFF; mem['h1F2D]=8'hFF; mem['h1F2E]=8'hFF; mem['h1F2F]=8'hFF;
    mem['h1F30]=8'hFF; mem['h1F31]=8'hFF; mem['h1F32]=8'hFF; mem['h1F33]=8'hFF;
    mem['h1F34]=8'hFF; mem['h1F35]=8'hFF; mem['h1F36]=8'hFF; mem['h1F37]=8'hFF;
    mem['h1F38]=8'hFF; mem['h1F39]=8'hFF; mem['h1F3A]=8'hFF; mem['h1F3B]=8'hFF;
    mem['h1F3C]=8'hFF; mem['h1F3D]=8'hFF; mem['h1F3E]=8'hFF; mem['h1F3F]=8'hFF;
    mem['h1F40]=8'hFF; mem['h1F41]=8'hFF; mem['h1F42]=8'hFF; mem['h1F43]=8'hFF;
    mem['h1F44]=8'hFF; mem['h1F45]=8'hFF; mem['h1F46]=8'hFF; mem['h1F47]=8'hFF;
    mem['h1F48]=8'hFF; mem['h1F49]=8'hFF; mem['h1F4A]=8'hFF; mem['h1F4B]=8'hFF;
    mem['h1F4C]=8'hFF; mem['h1F4D]=8'hFF; mem['h1F4E]=8'hFF; mem['h1F4F]=8'hFF;
    mem['h1F50]=8'hFF; mem['h1F51]=8'hFF; mem['h1F52]=8'hFF; mem['h1F53]=8'hFF;
    mem['h1F54]=8'hFF; mem['h1F55]=8'hFF; mem['h1F56]=8'hFF; mem['h1F57]=8'hFF;
    mem['h1F58]=8'hFF; mem['h1F59]=8'hFF; mem['h1F5A]=8'hFF; mem['h1F5B]=8'hFF;
    mem['h1F5C]=8'hFF; mem['h1F5D]=8'hFF; mem['h1F5E]=8'hFF; mem['h1F5F]=8'hFF;
    mem['h1F60]=8'hFF; mem['h1F61]=8'hFF; mem['h1F62]=8'hFF; mem['h1F63]=8'hFF;
    mem['h1F64]=8'hFF; mem['h1F65]=8'hFF; mem['h1F66]=8'hFF; mem['h1F67]=8'hFF;
    mem['h1F68]=8'hFF; mem['h1F69]=8'hFF; mem['h1F6A]=8'hFF; mem['h1F6B]=8'hFF;
    mem['h1F6C]=8'hFF; mem['h1F6D]=8'hFF; mem['h1F6E]=8'hFF; mem['h1F6F]=8'hFF;
    mem['h1F70]=8'hFF; mem['h1F71]=8'hFF; mem['h1F72]=8'hFF; mem['h1F73]=8'hFF;
    mem['h1F74]=8'hFF; mem['h1F75]=8'hFF; mem['h1F76]=8'hFF; mem['h1F77]=8'hFF;
    mem['h1F78]=8'hFF; mem['h1F79]=8'hFF; mem['h1F7A]=8'hFF; mem['h1F7B]=8'hFF;
    mem['h1F7C]=8'hFF; mem['h1F7D]=8'hFF; mem['h1F7E]=8'hFF; mem['h1F7F]=8'hFF;
    mem['h1F80]=8'hFF; mem['h1F81]=8'hFF; mem['h1F82]=8'hFF; mem['h1F83]=8'hFF;
    mem['h1F84]=8'hFF; mem['h1F85]=8'hFF; mem['h1F86]=8'hFF; mem['h1F87]=8'hFF;
    mem['h1F88]=8'hFF; mem['h1F89]=8'hFF; mem['h1F8A]=8'hFF; mem['h1F8B]=8'hFF;
    mem['h1F8C]=8'hFF; mem['h1F8D]=8'hFF; mem['h1F8E]=8'hFF; mem['h1F8F]=8'hFF;
    mem['h1F90]=8'hFF; mem['h1F91]=8'hFF; mem['h1F92]=8'hFF; mem['h1F93]=8'hFF;
    mem['h1F94]=8'hFF; mem['h1F95]=8'hFF; mem['h1F96]=8'hFF; mem['h1F97]=8'hFF;
    mem['h1F98]=8'hFF; mem['h1F99]=8'hFF; mem['h1F9A]=8'hFF; mem['h1F9B]=8'hFF;
    mem['h1F9C]=8'hFF; mem['h1F9D]=8'hFF; mem['h1F9E]=8'hFF; mem['h1F9F]=8'hFF;
    mem['h1FA0]=8'hFF; mem['h1FA1]=8'hFF; mem['h1FA2]=8'hFF; mem['h1FA3]=8'hFF;
    mem['h1FA4]=8'hFF; mem['h1FA5]=8'hFF; mem['h1FA6]=8'hFF; mem['h1FA7]=8'hFF;
    mem['h1FA8]=8'hFF; mem['h1FA9]=8'hFF; mem['h1FAA]=8'hFF; mem['h1FAB]=8'hFF;
    mem['h1FAC]=8'hFF; mem['h1FAD]=8'hFF; mem['h1FAE]=8'hFF; mem['h1FAF]=8'hFF;
    mem['h1FB0]=8'hFF; mem['h1FB1]=8'hFF; mem['h1FB2]=8'hFF; mem['h1FB3]=8'hFF;
    mem['h1FB4]=8'hFF; mem['h1FB5]=8'hFF; mem['h1FB6]=8'hFF; mem['h1FB7]=8'hFF;
    mem['h1FB8]=8'hFF; mem['h1FB9]=8'hFF; mem['h1FBA]=8'hFF; mem['h1FBB]=8'hFF;
    mem['h1FBC]=8'hFF; mem['h1FBD]=8'hFF; mem['h1FBE]=8'hFF; mem['h1FBF]=8'hFF;
    mem['h1FC0]=8'hFF; mem['h1FC1]=8'hFF; mem['h1FC2]=8'hFF; mem['h1FC3]=8'hFF;
    mem['h1FC4]=8'hFF; mem['h1FC5]=8'hFF; mem['h1FC6]=8'hFF; mem['h1FC7]=8'hFF;
    mem['h1FC8]=8'hFF; mem['h1FC9]=8'hFF; mem['h1FCA]=8'hFF; mem['h1FCB]=8'hFF;
    mem['h1FCC]=8'hFF; mem['h1FCD]=8'hFF; mem['h1FCE]=8'hFF; mem['h1FCF]=8'hFF;
    mem['h1FD0]=8'hFF; mem['h1FD1]=8'hFF; mem['h1FD2]=8'hFF; mem['h1FD3]=8'hFF;
    mem['h1FD4]=8'hFF; mem['h1FD5]=8'hFF; mem['h1FD6]=8'hFF; mem['h1FD7]=8'hFF;
    mem['h1FD8]=8'hFF; mem['h1FD9]=8'hFF; mem['h1FDA]=8'hFF; mem['h1FDB]=8'hFF;
    mem['h1FDC]=8'hFF; mem['h1FDD]=8'hFF; mem['h1FDE]=8'hFF; mem['h1FDF]=8'hFF;
    mem['h1FE0]=8'hFF; mem['h1FE1]=8'hFF; mem['h1FE2]=8'hFF; mem['h1FE3]=8'hFF;
    mem['h1FE4]=8'hFF; mem['h1FE5]=8'hFF; mem['h1FE6]=8'hFF; mem['h1FE7]=8'hFF;
    mem['h1FE8]=8'hFF; mem['h1FE9]=8'hFF; mem['h1FEA]=8'hFF; mem['h1FEB]=8'hFF;
    mem['h1FEC]=8'hFF; mem['h1FED]=8'hFF; mem['h1FEE]=8'hFF; mem['h1FEF]=8'hFF;
    mem['h1FF0]=8'hFF; mem['h1FF1]=8'hFF; mem['h1FF2]=8'hFF; mem['h1FF3]=8'hFF;
    mem['h1FF4]=8'hFF; mem['h1FF5]=8'hFF; mem['h1FF6]=8'hFF; mem['h1FF7]=8'hFF;
    mem['h1FF8]=8'hFF; mem['h1FF9]=8'hFF; mem['h1FFA]=8'hFF; mem['h1FFB]=8'hFF;
    mem['h1FFC]=8'hFF; mem['h1FFD]=8'hFF; mem['h1FFE]=8'hFF; mem['h1FFF]=8'hFF;
    mem['h2000]=8'h00; mem['h2001]=8'h00; mem['h2002]=8'h00; mem['h2003]=8'h00;
    mem['h2004]=8'h00; mem['h2005]=8'h00; mem['h2006]=8'h00; mem['h2007]=8'h00;
    mem['h2008]=8'h00; mem['h2009]=8'h00; mem['h200A]=8'h00; mem['h200B]=8'h00;
    mem['h200C]=8'h00; mem['h200D]=8'h00; mem['h200E]=8'h00; mem['h200F]=8'h00;
    mem['h2010]=8'h00; mem['h2011]=8'h00; mem['h2012]=8'h00; mem['h2013]=8'h00;
    mem['h2014]=8'h00; mem['h2015]=8'h00; mem['h2016]=8'h00; mem['h2017]=8'h00;
    mem['h2018]=8'h00; mem['h2019]=8'h00; mem['h201A]=8'h00; mem['h201B]=8'h00;
    mem['h201C]=8'h00; mem['h201D]=8'h00; mem['h201E]=8'h00; mem['h201F]=8'h00;
    mem['h2020]=8'h00; mem['h2021]=8'h00; mem['h2022]=8'h00; mem['h2023]=8'h00;
    mem['h2024]=8'h00; mem['h2025]=8'h00; mem['h2026]=8'h00; mem['h2027]=8'h00;
    mem['h2028]=8'h00; mem['h2029]=8'h00; mem['h202A]=8'h00; mem['h202B]=8'h00;
    mem['h202C]=8'h00; mem['h202D]=8'h00; mem['h202E]=8'h00; mem['h202F]=8'h00;
    mem['h2030]=8'h00; mem['h2031]=8'h00; mem['h2032]=8'h00; mem['h2033]=8'h00;
    mem['h2034]=8'h00; mem['h2035]=8'h00; mem['h2036]=8'h00; mem['h2037]=8'h00;
    mem['h2038]=8'h00; mem['h2039]=8'h00; mem['h203A]=8'h00; mem['h203B]=8'h00;
    mem['h203C]=8'h00; mem['h203D]=8'h00; mem['h203E]=8'h00; mem['h203F]=8'h00;
    mem['h2040]=8'h00; mem['h2041]=8'h00; mem['h2042]=8'h00; mem['h2043]=8'h00;
    mem['h2044]=8'h00; mem['h2045]=8'h00; mem['h2046]=8'h00; mem['h2047]=8'h00;
    mem['h2048]=8'h00; mem['h2049]=8'h00; mem['h204A]=8'h00; mem['h204B]=8'h00;
    mem['h204C]=8'h00; mem['h204D]=8'h00; mem['h204E]=8'h00; mem['h204F]=8'h00;
    mem['h2050]=8'h00; mem['h2051]=8'h00; mem['h2052]=8'h00; mem['h2053]=8'h00;
    mem['h2054]=8'h00; mem['h2055]=8'h00; mem['h2056]=8'h00; mem['h2057]=8'h00;
    mem['h2058]=8'h00; mem['h2059]=8'h00; mem['h205A]=8'h00; mem['h205B]=8'h00;
    mem['h205C]=8'h00; mem['h205D]=8'h00; mem['h205E]=8'h00; mem['h205F]=8'h00;
    mem['h2060]=8'h00; mem['h2061]=8'h00; mem['h2062]=8'h00; mem['h2063]=8'h00;
    mem['h2064]=8'h00; mem['h2065]=8'h00; mem['h2066]=8'h00; mem['h2067]=8'h00;
    mem['h2068]=8'h00; mem['h2069]=8'h00; mem['h206A]=8'h00; mem['h206B]=8'h00;
    mem['h206C]=8'h00; mem['h206D]=8'h00; mem['h206E]=8'h00; mem['h206F]=8'h00;
    mem['h2070]=8'h00; mem['h2071]=8'h00; mem['h2072]=8'h00; mem['h2073]=8'h00;
    mem['h2074]=8'h00; mem['h2075]=8'h00; mem['h2076]=8'h00; mem['h2077]=8'h00;
    mem['h2078]=8'h00; mem['h2079]=8'h00; mem['h207A]=8'h00; mem['h207B]=8'h00;
    mem['h207C]=8'h00; mem['h207D]=8'h00; mem['h207E]=8'h00; mem['h207F]=8'h00;
    mem['h2080]=8'h00; mem['h2081]=8'h00; mem['h2082]=8'h00; mem['h2083]=8'h00;
    mem['h2084]=8'h00; mem['h2085]=8'h00; mem['h2086]=8'h00; mem['h2087]=8'h00;
    mem['h2088]=8'h00; mem['h2089]=8'h00; mem['h208A]=8'h00; mem['h208B]=8'h00;
    mem['h208C]=8'h00; mem['h208D]=8'h00; mem['h208E]=8'h00; mem['h208F]=8'h00;
    mem['h2090]=8'h00; mem['h2091]=8'h00; mem['h2092]=8'h00; mem['h2093]=8'h00;
    mem['h2094]=8'h00; mem['h2095]=8'h00; mem['h2096]=8'h00; mem['h2097]=8'h00;
    mem['h2098]=8'h00; mem['h2099]=8'h00; mem['h209A]=8'h00; mem['h209B]=8'h00;
    mem['h209C]=8'h00; mem['h209D]=8'h00; mem['h209E]=8'h00; mem['h209F]=8'h00;
    mem['h20A0]=8'h00; mem['h20A1]=8'h00; mem['h20A2]=8'h00; mem['h20A3]=8'h00;
    mem['h20A4]=8'h00; mem['h20A5]=8'h00; mem['h20A6]=8'h00; mem['h20A7]=8'h00;
    mem['h20A8]=8'h00; mem['h20A9]=8'h00; mem['h20AA]=8'h00; mem['h20AB]=8'h00;
    mem['h20AC]=8'h00; mem['h20AD]=8'h00; mem['h20AE]=8'h00; mem['h20AF]=8'h00;
    mem['h20B0]=8'h00; mem['h20B1]=8'h00; mem['h20B2]=8'h00; mem['h20B3]=8'h00;
    mem['h20B4]=8'h00; mem['h20B5]=8'h00; mem['h20B6]=8'h00; mem['h20B7]=8'h00;
    mem['h20B8]=8'h00; mem['h20B9]=8'h00; mem['h20BA]=8'h00; mem['h20BB]=8'h00;
    mem['h20BC]=8'h00; mem['h20BD]=8'h00; mem['h20BE]=8'h00; mem['h20BF]=8'h00;
    mem['h20C0]=8'h00; mem['h20C1]=8'h00; mem['h20C2]=8'h00; mem['h20C3]=8'h00;
    mem['h20C4]=8'h00; mem['h20C5]=8'h00; mem['h20C6]=8'h00; mem['h20C7]=8'h00;
    mem['h20C8]=8'h00; mem['h20C9]=8'h00; mem['h20CA]=8'h00; mem['h20CB]=8'h00;
    mem['h20CC]=8'h00; mem['h20CD]=8'h00; mem['h20CE]=8'h00; mem['h20CF]=8'h00;
    mem['h20D0]=8'h00; mem['h20D1]=8'h00; mem['h20D2]=8'h00; mem['h20D3]=8'h00;
    mem['h20D4]=8'h00; mem['h20D5]=8'h00; mem['h20D6]=8'h00; mem['h20D7]=8'h00;
    mem['h20D8]=8'h00; mem['h20D9]=8'h00; mem['h20DA]=8'h00; mem['h20DB]=8'h00;
    mem['h20DC]=8'h00; mem['h20DD]=8'h00; mem['h20DE]=8'h00; mem['h20DF]=8'h00;
    mem['h20E0]=8'h00; mem['h20E1]=8'h00; mem['h20E2]=8'h00; mem['h20E3]=8'h00;
    mem['h20E4]=8'h00; mem['h20E5]=8'h00; mem['h20E6]=8'h00; mem['h20E7]=8'h00;
    mem['h20E8]=8'h00; mem['h20E9]=8'h00; mem['h20EA]=8'h00; mem['h20EB]=8'h00;
    mem['h20EC]=8'h00; mem['h20ED]=8'h00; mem['h20EE]=8'h00; mem['h20EF]=8'h00;
    mem['h20F0]=8'h00; mem['h20F1]=8'h00; mem['h20F2]=8'h00; mem['h20F3]=8'h00;
    mem['h20F4]=8'h00; mem['h20F5]=8'h00; mem['h20F6]=8'h00; mem['h20F7]=8'h00;
    mem['h20F8]=8'h00; mem['h20F9]=8'h00; mem['h20FA]=8'h00; mem['h20FB]=8'h00;
    mem['h20FC]=8'h00; mem['h20FD]=8'h00; mem['h20FE]=8'h00; mem['h20FF]=8'h00;
    mem['h2100]=8'h00; mem['h2101]=8'h00; mem['h2102]=8'h00; mem['h2103]=8'h00;
    mem['h2104]=8'h00; mem['h2105]=8'h00; mem['h2106]=8'h00; mem['h2107]=8'h00;
    mem['h2108]=8'h00; mem['h2109]=8'h00; mem['h210A]=8'h00; mem['h210B]=8'h00;
    mem['h210C]=8'h00; mem['h210D]=8'h00; mem['h210E]=8'h00; mem['h210F]=8'h00;
    mem['h2110]=8'h00; mem['h2111]=8'h00; mem['h2112]=8'h00; mem['h2113]=8'h00;
    mem['h2114]=8'h00; mem['h2115]=8'h00; mem['h2116]=8'h00; mem['h2117]=8'h00;
    mem['h2118]=8'h00; mem['h2119]=8'h00; mem['h211A]=8'h00; mem['h211B]=8'h00;
    mem['h211C]=8'h00; mem['h211D]=8'h00; mem['h211E]=8'h00; mem['h211F]=8'h00;
    mem['h2120]=8'h00; mem['h2121]=8'h00; mem['h2122]=8'h00; mem['h2123]=8'h00;
    mem['h2124]=8'h00; mem['h2125]=8'h00; mem['h2126]=8'h00; mem['h2127]=8'h00;
    mem['h2128]=8'h00; mem['h2129]=8'h00; mem['h212A]=8'h00; mem['h212B]=8'h00;
    mem['h212C]=8'h00; mem['h212D]=8'h00; mem['h212E]=8'h00; mem['h212F]=8'h00;
    mem['h2130]=8'h00; mem['h2131]=8'h00; mem['h2132]=8'h00; mem['h2133]=8'h00;
    mem['h2134]=8'h00; mem['h2135]=8'h00; mem['h2136]=8'h00; mem['h2137]=8'h00;
    mem['h2138]=8'h00; mem['h2139]=8'h00; mem['h213A]=8'h00; mem['h213B]=8'h00;
    mem['h213C]=8'h00; mem['h213D]=8'h00; mem['h213E]=8'h00; mem['h213F]=8'h00;
    mem['h2140]=8'h00; mem['h2141]=8'h00; mem['h2142]=8'h00; mem['h2143]=8'h00;
    mem['h2144]=8'h00; mem['h2145]=8'h00; mem['h2146]=8'h00; mem['h2147]=8'h00;
    mem['h2148]=8'h00; mem['h2149]=8'h00; mem['h214A]=8'h00; mem['h214B]=8'h00;
    mem['h214C]=8'h00; mem['h214D]=8'h00; mem['h214E]=8'h00; mem['h214F]=8'h00;
    mem['h2150]=8'h00; mem['h2151]=8'h00; mem['h2152]=8'h00; mem['h2153]=8'h00;
    mem['h2154]=8'h00; mem['h2155]=8'h00; mem['h2156]=8'h00; mem['h2157]=8'h00;
    mem['h2158]=8'h00; mem['h2159]=8'h00; mem['h215A]=8'h00; mem['h215B]=8'h00;
    mem['h215C]=8'h00; mem['h215D]=8'h00; mem['h215E]=8'h00; mem['h215F]=8'h00;
    mem['h2160]=8'h00; mem['h2161]=8'h00; mem['h2162]=8'h00; mem['h2163]=8'h00;
    mem['h2164]=8'h00; mem['h2165]=8'h00; mem['h2166]=8'h00; mem['h2167]=8'h00;
    mem['h2168]=8'h00; mem['h2169]=8'h00; mem['h216A]=8'h00; mem['h216B]=8'h00;
    mem['h216C]=8'h00; mem['h216D]=8'h00; mem['h216E]=8'h00; mem['h216F]=8'h00;
    mem['h2170]=8'h00; mem['h2171]=8'h00; mem['h2172]=8'h00; mem['h2173]=8'h00;
    mem['h2174]=8'h00; mem['h2175]=8'h00; mem['h2176]=8'h00; mem['h2177]=8'h00;
    mem['h2178]=8'h00; mem['h2179]=8'h00; mem['h217A]=8'h00; mem['h217B]=8'h00;
    mem['h217C]=8'h00; mem['h217D]=8'h00; mem['h217E]=8'h00; mem['h217F]=8'h00;
    mem['h2180]=8'h00; mem['h2181]=8'h00; mem['h2182]=8'h00; mem['h2183]=8'h00;
    mem['h2184]=8'h00; mem['h2185]=8'h00; mem['h2186]=8'h00; mem['h2187]=8'h00;
    mem['h2188]=8'h00; mem['h2189]=8'h00; mem['h218A]=8'h00; mem['h218B]=8'h00;
    mem['h218C]=8'h00; mem['h218D]=8'h00; mem['h218E]=8'h00; mem['h218F]=8'h00;
    mem['h2190]=8'h00; mem['h2191]=8'h00; mem['h2192]=8'h00; mem['h2193]=8'h00;
    mem['h2194]=8'h00; mem['h2195]=8'h00; mem['h2196]=8'h00; mem['h2197]=8'h00;
    mem['h2198]=8'h00; mem['h2199]=8'h00; mem['h219A]=8'h00; mem['h219B]=8'h00;
    mem['h219C]=8'h00; mem['h219D]=8'h00; mem['h219E]=8'h00; mem['h219F]=8'h00;
    mem['h21A0]=8'h00; mem['h21A1]=8'h00; mem['h21A2]=8'h00; mem['h21A3]=8'h00;
    mem['h21A4]=8'h00; mem['h21A5]=8'h00; mem['h21A6]=8'h00; mem['h21A7]=8'h00;
    mem['h21A8]=8'h00; mem['h21A9]=8'h00; mem['h21AA]=8'h00; mem['h21AB]=8'h00;
    mem['h21AC]=8'h00; mem['h21AD]=8'h00; mem['h21AE]=8'h00; mem['h21AF]=8'h00;
    mem['h21B0]=8'h00; mem['h21B1]=8'h00; mem['h21B2]=8'h00; mem['h21B3]=8'h00;
    mem['h21B4]=8'h00; mem['h21B5]=8'h00; mem['h21B6]=8'h00; mem['h21B7]=8'h00;
    mem['h21B8]=8'h00; mem['h21B9]=8'h00; mem['h21BA]=8'h00; mem['h21BB]=8'h00;
    mem['h21BC]=8'h00; mem['h21BD]=8'h00; mem['h21BE]=8'h00; mem['h21BF]=8'h00;
    mem['h21C0]=8'h00; mem['h21C1]=8'h00; mem['h21C2]=8'h00; mem['h21C3]=8'h00;
    mem['h21C4]=8'h00; mem['h21C5]=8'h00; mem['h21C6]=8'h00; mem['h21C7]=8'h00;
    mem['h21C8]=8'h00; mem['h21C9]=8'h00; mem['h21CA]=8'h00; mem['h21CB]=8'h00;
    mem['h21CC]=8'h00; mem['h21CD]=8'h00; mem['h21CE]=8'h00; mem['h21CF]=8'h00;
    mem['h21D0]=8'h00; mem['h21D1]=8'h00; mem['h21D2]=8'h00; mem['h21D3]=8'h00;
    mem['h21D4]=8'h00; mem['h21D5]=8'h00; mem['h21D6]=8'h00; mem['h21D7]=8'h00;
    mem['h21D8]=8'h00; mem['h21D9]=8'h00; mem['h21DA]=8'h00; mem['h21DB]=8'h00;
    mem['h21DC]=8'h00; mem['h21DD]=8'h00; mem['h21DE]=8'h00; mem['h21DF]=8'h00;
    mem['h21E0]=8'h00; mem['h21E1]=8'h00; mem['h21E2]=8'h00; mem['h21E3]=8'h00;
    mem['h21E4]=8'h00; mem['h21E5]=8'h00; mem['h21E6]=8'h00; mem['h21E7]=8'h00;
    mem['h21E8]=8'h00; mem['h21E9]=8'h00; mem['h21EA]=8'h00; mem['h21EB]=8'h00;
    mem['h21EC]=8'h00; mem['h21ED]=8'h00; mem['h21EE]=8'h00; mem['h21EF]=8'h00;
    mem['h21F0]=8'h00; mem['h21F1]=8'h00; mem['h21F2]=8'h00; mem['h21F3]=8'h00;
    mem['h21F4]=8'h00; mem['h21F5]=8'h00; mem['h21F6]=8'h00; mem['h21F7]=8'h00;
    mem['h21F8]=8'h00; mem['h21F9]=8'h00; mem['h21FA]=8'h00; mem['h21FB]=8'h00;
    mem['h21FC]=8'h00; mem['h21FD]=8'h00; mem['h21FE]=8'h00; mem['h21FF]=8'h00;
    mem['h2200]=8'h00; mem['h2201]=8'h00; mem['h2202]=8'h00; mem['h2203]=8'h00;
    mem['h2204]=8'h00; mem['h2205]=8'h00; mem['h2206]=8'h00; mem['h2207]=8'h00;
    mem['h2208]=8'h00; mem['h2209]=8'h00; mem['h220A]=8'h00; mem['h220B]=8'h00;
    mem['h220C]=8'h00; mem['h220D]=8'h00; mem['h220E]=8'h00; mem['h220F]=8'h00;
    mem['h2210]=8'h00; mem['h2211]=8'h00; mem['h2212]=8'h00; mem['h2213]=8'h00;
    mem['h2214]=8'h00; mem['h2215]=8'h00; mem['h2216]=8'h00; mem['h2217]=8'h00;
    mem['h2218]=8'h00; mem['h2219]=8'h00; mem['h221A]=8'h00; mem['h221B]=8'h00;
    mem['h221C]=8'h00; mem['h221D]=8'h00; mem['h221E]=8'h00; mem['h221F]=8'h00;
    mem['h2220]=8'h00; mem['h2221]=8'h00; mem['h2222]=8'h00; mem['h2223]=8'h00;
    mem['h2224]=8'h00; mem['h2225]=8'h00; mem['h2226]=8'h00; mem['h2227]=8'h00;
    mem['h2228]=8'h00; mem['h2229]=8'h00; mem['h222A]=8'h00; mem['h222B]=8'h00;
    mem['h222C]=8'h00; mem['h222D]=8'h00; mem['h222E]=8'h00; mem['h222F]=8'h00;
    mem['h2230]=8'h00; mem['h2231]=8'h00; mem['h2232]=8'h00; mem['h2233]=8'h00;
    mem['h2234]=8'h00; mem['h2235]=8'h00; mem['h2236]=8'h00; mem['h2237]=8'h00;
    mem['h2238]=8'h00; mem['h2239]=8'h00; mem['h223A]=8'h00; mem['h223B]=8'h00;
    mem['h223C]=8'h00; mem['h223D]=8'h00; mem['h223E]=8'h00; mem['h223F]=8'h00;
    mem['h2240]=8'h00; mem['h2241]=8'h00; mem['h2242]=8'h00; mem['h2243]=8'h00;
    mem['h2244]=8'h00; mem['h2245]=8'h00; mem['h2246]=8'h00; mem['h2247]=8'h00;
    mem['h2248]=8'h00; mem['h2249]=8'h00; mem['h224A]=8'h00; mem['h224B]=8'h00;
    mem['h224C]=8'h00; mem['h224D]=8'h00; mem['h224E]=8'h00; mem['h224F]=8'h00;
    mem['h2250]=8'h00; mem['h2251]=8'h00; mem['h2252]=8'h00; mem['h2253]=8'h00;
    mem['h2254]=8'h00; mem['h2255]=8'h00; mem['h2256]=8'h00; mem['h2257]=8'h00;
    mem['h2258]=8'h00; mem['h2259]=8'h00; mem['h225A]=8'h00; mem['h225B]=8'h00;
    mem['h225C]=8'h00; mem['h225D]=8'h00; mem['h225E]=8'h00; mem['h225F]=8'h00;
    mem['h2260]=8'h00; mem['h2261]=8'h00; mem['h2262]=8'h00; mem['h2263]=8'h00;
    mem['h2264]=8'h00; mem['h2265]=8'h00; mem['h2266]=8'h00; mem['h2267]=8'h00;
    mem['h2268]=8'h00; mem['h2269]=8'h00; mem['h226A]=8'h00; mem['h226B]=8'h00;
    mem['h226C]=8'h00; mem['h226D]=8'h00; mem['h226E]=8'h00; mem['h226F]=8'h00;
    mem['h2270]=8'h00; mem['h2271]=8'h00; mem['h2272]=8'h00; mem['h2273]=8'h00;
    mem['h2274]=8'h00; mem['h2275]=8'h00; mem['h2276]=8'h00; mem['h2277]=8'h00;
    mem['h2278]=8'h00; mem['h2279]=8'h00; mem['h227A]=8'h00; mem['h227B]=8'h00;
    mem['h227C]=8'h00; mem['h227D]=8'h00; mem['h227E]=8'h00; mem['h227F]=8'h00;
    mem['h2280]=8'h00; mem['h2281]=8'h00; mem['h2282]=8'h00; mem['h2283]=8'h00;
    mem['h2284]=8'h00; mem['h2285]=8'h00; mem['h2286]=8'h00; mem['h2287]=8'h00;
    mem['h2288]=8'h00; mem['h2289]=8'h00; mem['h228A]=8'h00; mem['h228B]=8'h00;
    mem['h228C]=8'h00; mem['h228D]=8'h00; mem['h228E]=8'h00; mem['h228F]=8'h00;
    mem['h2290]=8'h00; mem['h2291]=8'h00; mem['h2292]=8'h00; mem['h2293]=8'h00;
    mem['h2294]=8'h00; mem['h2295]=8'h00; mem['h2296]=8'h00; mem['h2297]=8'h00;
    mem['h2298]=8'h00; mem['h2299]=8'h00; mem['h229A]=8'h00; mem['h229B]=8'h00;
    mem['h229C]=8'h00; mem['h229D]=8'h00; mem['h229E]=8'h00; mem['h229F]=8'h00;
    mem['h22A0]=8'h00; mem['h22A1]=8'h00; mem['h22A2]=8'h00; mem['h22A3]=8'h00;
    mem['h22A4]=8'h00; mem['h22A5]=8'h00; mem['h22A6]=8'h00; mem['h22A7]=8'h00;
    mem['h22A8]=8'h00; mem['h22A9]=8'h00; mem['h22AA]=8'h00; mem['h22AB]=8'h00;
    mem['h22AC]=8'h00; mem['h22AD]=8'h00; mem['h22AE]=8'h00; mem['h22AF]=8'h00;
    mem['h22B0]=8'h00; mem['h22B1]=8'h00; mem['h22B2]=8'h00; mem['h22B3]=8'h00;
    mem['h22B4]=8'h00; mem['h22B5]=8'h00; mem['h22B6]=8'h00; mem['h22B7]=8'h00;
    mem['h22B8]=8'h00; mem['h22B9]=8'h00; mem['h22BA]=8'h00; mem['h22BB]=8'h00;
    mem['h22BC]=8'h00; mem['h22BD]=8'h00; mem['h22BE]=8'h00; mem['h22BF]=8'h00;
    mem['h22C0]=8'h00; mem['h22C1]=8'h00; mem['h22C2]=8'h00; mem['h22C3]=8'h00;
    mem['h22C4]=8'h00; mem['h22C5]=8'h00; mem['h22C6]=8'h00; mem['h22C7]=8'h00;
    mem['h22C8]=8'h00; mem['h22C9]=8'h00; mem['h22CA]=8'h00; mem['h22CB]=8'h00;
    mem['h22CC]=8'h00; mem['h22CD]=8'h00; mem['h22CE]=8'h00; mem['h22CF]=8'h00;
    mem['h22D0]=8'h00; mem['h22D1]=8'h00; mem['h22D2]=8'h00; mem['h22D3]=8'h00;
    mem['h22D4]=8'h00; mem['h22D5]=8'h00; mem['h22D6]=8'h00; mem['h22D7]=8'h00;
    mem['h22D8]=8'h00; mem['h22D9]=8'h00; mem['h22DA]=8'h00; mem['h22DB]=8'h00;
    mem['h22DC]=8'h00; mem['h22DD]=8'h00; mem['h22DE]=8'h00; mem['h22DF]=8'h00;
    mem['h22E0]=8'h00; mem['h22E1]=8'h00; mem['h22E2]=8'h00; mem['h22E3]=8'h00;
    mem['h22E4]=8'h00; mem['h22E5]=8'h00; mem['h22E6]=8'h00; mem['h22E7]=8'h00;
    mem['h22E8]=8'h00; mem['h22E9]=8'h00; mem['h22EA]=8'h00; mem['h22EB]=8'h00;
    mem['h22EC]=8'h00; mem['h22ED]=8'h00; mem['h22EE]=8'h00; mem['h22EF]=8'h00;
    mem['h22F0]=8'h00; mem['h22F1]=8'h00; mem['h22F2]=8'h00; mem['h22F3]=8'h00;
    mem['h22F4]=8'h00; mem['h22F5]=8'h00; mem['h22F6]=8'h00; mem['h22F7]=8'h00;
    mem['h22F8]=8'h00; mem['h22F9]=8'h00; mem['h22FA]=8'h00; mem['h22FB]=8'h00;
    mem['h22FC]=8'h00; mem['h22FD]=8'h00; mem['h22FE]=8'h00; mem['h22FF]=8'h00;
    mem['h2300]=8'h00; mem['h2301]=8'h00; mem['h2302]=8'h00; mem['h2303]=8'h00;
    mem['h2304]=8'h00; mem['h2305]=8'h00; mem['h2306]=8'h00; mem['h2307]=8'h00;
    mem['h2308]=8'h00; mem['h2309]=8'h00; mem['h230A]=8'h00; mem['h230B]=8'h00;
    mem['h230C]=8'h00; mem['h230D]=8'h00; mem['h230E]=8'h00; mem['h230F]=8'h00;
    mem['h2310]=8'h00; mem['h2311]=8'h00; mem['h2312]=8'h00; mem['h2313]=8'h00;
    mem['h2314]=8'h00; mem['h2315]=8'h00; mem['h2316]=8'h00; mem['h2317]=8'h00;
    mem['h2318]=8'h00; mem['h2319]=8'h00; mem['h231A]=8'h00; mem['h231B]=8'h00;
    mem['h231C]=8'h00; mem['h231D]=8'h00; mem['h231E]=8'h00; mem['h231F]=8'h00;
    mem['h2320]=8'h00; mem['h2321]=8'h00; mem['h2322]=8'h00; mem['h2323]=8'h00;
    mem['h2324]=8'h00; mem['h2325]=8'h00; mem['h2326]=8'h00; mem['h2327]=8'h00;
    mem['h2328]=8'h00; mem['h2329]=8'h00; mem['h232A]=8'h00; mem['h232B]=8'h00;
    mem['h232C]=8'h00; mem['h232D]=8'h00; mem['h232E]=8'h00; mem['h232F]=8'h00;
    mem['h2330]=8'h00; mem['h2331]=8'h00; mem['h2332]=8'h00; mem['h2333]=8'h00;
    mem['h2334]=8'h00; mem['h2335]=8'h00; mem['h2336]=8'h00; mem['h2337]=8'h00;
    mem['h2338]=8'h00; mem['h2339]=8'h00; mem['h233A]=8'h00; mem['h233B]=8'h00;
    mem['h233C]=8'h00; mem['h233D]=8'h00; mem['h233E]=8'h00; mem['h233F]=8'h00;
    mem['h2340]=8'h00; mem['h2341]=8'h00; mem['h2342]=8'h00; mem['h2343]=8'h00;
    mem['h2344]=8'h00; mem['h2345]=8'h00; mem['h2346]=8'h00; mem['h2347]=8'h00;
    mem['h2348]=8'h00; mem['h2349]=8'h00; mem['h234A]=8'h00; mem['h234B]=8'h00;
    mem['h234C]=8'h00; mem['h234D]=8'h00; mem['h234E]=8'h00; mem['h234F]=8'h00;
    mem['h2350]=8'h00; mem['h2351]=8'h00; mem['h2352]=8'h00; mem['h2353]=8'h00;
    mem['h2354]=8'h00; mem['h2355]=8'h00; mem['h2356]=8'h00; mem['h2357]=8'h00;
    mem['h2358]=8'h00; mem['h2359]=8'h00; mem['h235A]=8'h00; mem['h235B]=8'h00;
    mem['h235C]=8'h00; mem['h235D]=8'h00; mem['h235E]=8'h00; mem['h235F]=8'h00;
    mem['h2360]=8'h00; mem['h2361]=8'h00; mem['h2362]=8'h00; mem['h2363]=8'h00;
    mem['h2364]=8'h00; mem['h2365]=8'h00; mem['h2366]=8'h00; mem['h2367]=8'h00;
    mem['h2368]=8'h00; mem['h2369]=8'h00; mem['h236A]=8'h00; mem['h236B]=8'h00;
    mem['h236C]=8'h00; mem['h236D]=8'h00; mem['h236E]=8'h00; mem['h236F]=8'h00;
    mem['h2370]=8'h00; mem['h2371]=8'h00; mem['h2372]=8'h00; mem['h2373]=8'h00;
    mem['h2374]=8'h00; mem['h2375]=8'h00; mem['h2376]=8'h00; mem['h2377]=8'h00;
    mem['h2378]=8'h00; mem['h2379]=8'h00; mem['h237A]=8'h00; mem['h237B]=8'h00;
    mem['h237C]=8'h00; mem['h237D]=8'h00; mem['h237E]=8'h00; mem['h237F]=8'h00;
    mem['h2380]=8'h00; mem['h2381]=8'h00; mem['h2382]=8'h00; mem['h2383]=8'h00;
    mem['h2384]=8'h00; mem['h2385]=8'h00; mem['h2386]=8'h00; mem['h2387]=8'h00;
    mem['h2388]=8'h00; mem['h2389]=8'h00; mem['h238A]=8'h00; mem['h238B]=8'h00;
    mem['h238C]=8'h00; mem['h238D]=8'h00; mem['h238E]=8'h00; mem['h238F]=8'h00;
    mem['h2390]=8'h00; mem['h2391]=8'h00; mem['h2392]=8'h00; mem['h2393]=8'h00;
    mem['h2394]=8'h00; mem['h2395]=8'h00; mem['h2396]=8'h00; mem['h2397]=8'h00;
    mem['h2398]=8'h00; mem['h2399]=8'h00; mem['h239A]=8'h00; mem['h239B]=8'h00;
    mem['h239C]=8'h00; mem['h239D]=8'h00; mem['h239E]=8'h00; mem['h239F]=8'h00;
    mem['h23A0]=8'h00; mem['h23A1]=8'h00; mem['h23A2]=8'h00; mem['h23A3]=8'h00;
    mem['h23A4]=8'h00; mem['h23A5]=8'h00; mem['h23A6]=8'h00; mem['h23A7]=8'h00;
    mem['h23A8]=8'h00; mem['h23A9]=8'h00; mem['h23AA]=8'h00; mem['h23AB]=8'h00;
    mem['h23AC]=8'h00; mem['h23AD]=8'h00; mem['h23AE]=8'h00; mem['h23AF]=8'h00;
    mem['h23B0]=8'h00; mem['h23B1]=8'h00; mem['h23B2]=8'h00; mem['h23B3]=8'h00;
    mem['h23B4]=8'h00; mem['h23B5]=8'h00; mem['h23B6]=8'h00; mem['h23B7]=8'h00;
    mem['h23B8]=8'h00; mem['h23B9]=8'h00; mem['h23BA]=8'h00; mem['h23BB]=8'h00;
    mem['h23BC]=8'h00; mem['h23BD]=8'h00; mem['h23BE]=8'h00; mem['h23BF]=8'h00;
    mem['h23C0]=8'h00; mem['h23C1]=8'h00; mem['h23C2]=8'h00; mem['h23C3]=8'h00;
    mem['h23C4]=8'h00; mem['h23C5]=8'h00; mem['h23C6]=8'h00; mem['h23C7]=8'h00;
    mem['h23C8]=8'h00; mem['h23C9]=8'h00; mem['h23CA]=8'h00; mem['h23CB]=8'h00;
    mem['h23CC]=8'h00; mem['h23CD]=8'h00; mem['h23CE]=8'h00; mem['h23CF]=8'h00;
    mem['h23D0]=8'h00; mem['h23D1]=8'h00; mem['h23D2]=8'h00; mem['h23D3]=8'h00;
    mem['h23D4]=8'h00; mem['h23D5]=8'h00; mem['h23D6]=8'h00; mem['h23D7]=8'h00;
    mem['h23D8]=8'h00; mem['h23D9]=8'h00; mem['h23DA]=8'h00; mem['h23DB]=8'h00;
    mem['h23DC]=8'h00; mem['h23DD]=8'h00; mem['h23DE]=8'h00; mem['h23DF]=8'h00;
    mem['h23E0]=8'h00; mem['h23E1]=8'h00; mem['h23E2]=8'h00; mem['h23E3]=8'h00;
    mem['h23E4]=8'h00; mem['h23E5]=8'h00; mem['h23E6]=8'h00; mem['h23E7]=8'h00;
    mem['h23E8]=8'h00; mem['h23E9]=8'h00; mem['h23EA]=8'h00; mem['h23EB]=8'h00;
    mem['h23EC]=8'h00; mem['h23ED]=8'h00; mem['h23EE]=8'h00; mem['h23EF]=8'h00;
    mem['h23F0]=8'h00; mem['h23F1]=8'h00; mem['h23F2]=8'h00; mem['h23F3]=8'h00;
    mem['h23F4]=8'h00; mem['h23F5]=8'h00; mem['h23F6]=8'h00; mem['h23F7]=8'h00;
    mem['h23F8]=8'h00; mem['h23F9]=8'h00; mem['h23FA]=8'h00; mem['h23FB]=8'h00;
    mem['h23FC]=8'h00; mem['h23FD]=8'h00; mem['h23FE]=8'h00; mem['h23FF]=8'h00;
    mem['h2400]=8'h00; mem['h2401]=8'h00; mem['h2402]=8'h00; mem['h2403]=8'h00;
    mem['h2404]=8'h00; mem['h2405]=8'h00; mem['h2406]=8'h00; mem['h2407]=8'h00;
    mem['h2408]=8'h00; mem['h2409]=8'h00; mem['h240A]=8'h00; mem['h240B]=8'h00;
    mem['h240C]=8'h00; mem['h240D]=8'h00; mem['h240E]=8'h00; mem['h240F]=8'h00;
    mem['h2410]=8'h00; mem['h2411]=8'h00; mem['h2412]=8'h00; mem['h2413]=8'h00;
    mem['h2414]=8'h00; mem['h2415]=8'h00; mem['h2416]=8'h00; mem['h2417]=8'h00;
    mem['h2418]=8'h00; mem['h2419]=8'h00; mem['h241A]=8'h00; mem['h241B]=8'h00;
    mem['h241C]=8'h00; mem['h241D]=8'h00; mem['h241E]=8'h00; mem['h241F]=8'h00;
    mem['h2420]=8'h00; mem['h2421]=8'h00; mem['h2422]=8'h00; mem['h2423]=8'h00;
    mem['h2424]=8'h00; mem['h2425]=8'h00; mem['h2426]=8'h00; mem['h2427]=8'h00;
    mem['h2428]=8'h00; mem['h2429]=8'h00; mem['h242A]=8'h00; mem['h242B]=8'h00;
    mem['h242C]=8'h00; mem['h242D]=8'h00; mem['h242E]=8'h00; mem['h242F]=8'h00;
    mem['h2430]=8'h00; mem['h2431]=8'h00; mem['h2432]=8'h00; mem['h2433]=8'h00;
    mem['h2434]=8'h00; mem['h2435]=8'h00; mem['h2436]=8'h00; mem['h2437]=8'h00;
    mem['h2438]=8'h00; mem['h2439]=8'h00; mem['h243A]=8'h00; mem['h243B]=8'h00;
    mem['h243C]=8'h00; mem['h243D]=8'h00; mem['h243E]=8'h00; mem['h243F]=8'h00;
    mem['h2440]=8'h00; mem['h2441]=8'h00; mem['h2442]=8'h00; mem['h2443]=8'h00;
    mem['h2444]=8'h00; mem['h2445]=8'h00; mem['h2446]=8'h00; mem['h2447]=8'h00;
    mem['h2448]=8'h00; mem['h2449]=8'h00; mem['h244A]=8'h00; mem['h244B]=8'h00;
    mem['h244C]=8'h00; mem['h244D]=8'h00; mem['h244E]=8'h00; mem['h244F]=8'h00;
    mem['h2450]=8'h00; mem['h2451]=8'h00; mem['h2452]=8'h00; mem['h2453]=8'h00;
    mem['h2454]=8'h00; mem['h2455]=8'h00; mem['h2456]=8'h00; mem['h2457]=8'h00;
    mem['h2458]=8'h00; mem['h2459]=8'h00; mem['h245A]=8'h00; mem['h245B]=8'h00;
    mem['h245C]=8'h00; mem['h245D]=8'h00; mem['h245E]=8'h00; mem['h245F]=8'h00;
    mem['h2460]=8'h00; mem['h2461]=8'h00; mem['h2462]=8'h00; mem['h2463]=8'h00;
    mem['h2464]=8'h00; mem['h2465]=8'h00; mem['h2466]=8'h00; mem['h2467]=8'h00;
    mem['h2468]=8'h00; mem['h2469]=8'h00; mem['h246A]=8'h00; mem['h246B]=8'h00;
    mem['h246C]=8'h00; mem['h246D]=8'h00; mem['h246E]=8'h00; mem['h246F]=8'h00;
    mem['h2470]=8'h00; mem['h2471]=8'h00; mem['h2472]=8'h00; mem['h2473]=8'h00;
    mem['h2474]=8'h00; mem['h2475]=8'h00; mem['h2476]=8'h00; mem['h2477]=8'h00;
    mem['h2478]=8'h00; mem['h2479]=8'h00; mem['h247A]=8'h00; mem['h247B]=8'h00;
    mem['h247C]=8'h00; mem['h247D]=8'h00; mem['h247E]=8'h00; mem['h247F]=8'h00;
    mem['h2480]=8'h00; mem['h2481]=8'h00; mem['h2482]=8'h00; mem['h2483]=8'h00;
    mem['h2484]=8'h00; mem['h2485]=8'h00; mem['h2486]=8'h00; mem['h2487]=8'h00;
    mem['h2488]=8'h00; mem['h2489]=8'h00; mem['h248A]=8'h00; mem['h248B]=8'h00;
    mem['h248C]=8'h00; mem['h248D]=8'h00; mem['h248E]=8'h00; mem['h248F]=8'h00;
    mem['h2490]=8'h00; mem['h2491]=8'h00; mem['h2492]=8'h00; mem['h2493]=8'h00;
    mem['h2494]=8'h00; mem['h2495]=8'h00; mem['h2496]=8'h00; mem['h2497]=8'h00;
    mem['h2498]=8'h00; mem['h2499]=8'h00; mem['h249A]=8'h00; mem['h249B]=8'h00;
    mem['h249C]=8'h00; mem['h249D]=8'h00; mem['h249E]=8'h00; mem['h249F]=8'h00;
    mem['h24A0]=8'h00; mem['h24A1]=8'h00; mem['h24A2]=8'h00; mem['h24A3]=8'h00;
    mem['h24A4]=8'h00; mem['h24A5]=8'h00; mem['h24A6]=8'h00; mem['h24A7]=8'h00;
    mem['h24A8]=8'h00; mem['h24A9]=8'h00; mem['h24AA]=8'h00; mem['h24AB]=8'h00;
    mem['h24AC]=8'h00; mem['h24AD]=8'h00; mem['h24AE]=8'h00; mem['h24AF]=8'h00;
    mem['h24B0]=8'h00; mem['h24B1]=8'h00; mem['h24B2]=8'h00; mem['h24B3]=8'h00;
    mem['h24B4]=8'h00; mem['h24B5]=8'h00; mem['h24B6]=8'h00; mem['h24B7]=8'h00;
    mem['h24B8]=8'h00; mem['h24B9]=8'h00; mem['h24BA]=8'h00; mem['h24BB]=8'h00;
    mem['h24BC]=8'h00; mem['h24BD]=8'h00; mem['h24BE]=8'h00; mem['h24BF]=8'h00;
    mem['h24C0]=8'h00; mem['h24C1]=8'h00; mem['h24C2]=8'h00; mem['h24C3]=8'h00;
    mem['h24C4]=8'h00; mem['h24C5]=8'h00; mem['h24C6]=8'h00; mem['h24C7]=8'h00;
    mem['h24C8]=8'h00; mem['h24C9]=8'h00; mem['h24CA]=8'h00; mem['h24CB]=8'h00;
    mem['h24CC]=8'h00; mem['h24CD]=8'h00; mem['h24CE]=8'h00; mem['h24CF]=8'h00;
    mem['h24D0]=8'h00; mem['h24D1]=8'h00; mem['h24D2]=8'h00; mem['h24D3]=8'h00;
    mem['h24D4]=8'h00; mem['h24D5]=8'h00; mem['h24D6]=8'h00; mem['h24D7]=8'h00;
    mem['h24D8]=8'h00; mem['h24D9]=8'h00; mem['h24DA]=8'h00; mem['h24DB]=8'h00;
    mem['h24DC]=8'h00; mem['h24DD]=8'h00; mem['h24DE]=8'h00; mem['h24DF]=8'h00;
    mem['h24E0]=8'h00; mem['h24E1]=8'h00; mem['h24E2]=8'h00; mem['h24E3]=8'h00;
    mem['h24E4]=8'h00; mem['h24E5]=8'h00; mem['h24E6]=8'h00; mem['h24E7]=8'h00;
    mem['h24E8]=8'h00; mem['h24E9]=8'h00; mem['h24EA]=8'h00; mem['h24EB]=8'h00;
    mem['h24EC]=8'h00; mem['h24ED]=8'h00; mem['h24EE]=8'h00; mem['h24EF]=8'h00;
    mem['h24F0]=8'h00; mem['h24F1]=8'h00; mem['h24F2]=8'h00; mem['h24F3]=8'h00;
    mem['h24F4]=8'h00; mem['h24F5]=8'h00; mem['h24F6]=8'h00; mem['h24F7]=8'h00;
    mem['h24F8]=8'h00; mem['h24F9]=8'h00; mem['h24FA]=8'h00; mem['h24FB]=8'h00;
    mem['h24FC]=8'h00; mem['h24FD]=8'h00; mem['h24FE]=8'h00; mem['h24FF]=8'h00;
    mem['h2500]=8'h00; mem['h2501]=8'h00; mem['h2502]=8'h00; mem['h2503]=8'h00;
    mem['h2504]=8'h00; mem['h2505]=8'h00; mem['h2506]=8'h00; mem['h2507]=8'h00;
    mem['h2508]=8'h00; mem['h2509]=8'h00; mem['h250A]=8'h00; mem['h250B]=8'h00;
    mem['h250C]=8'h00; mem['h250D]=8'h00; mem['h250E]=8'h00; mem['h250F]=8'h00;
    mem['h2510]=8'h00; mem['h2511]=8'h00; mem['h2512]=8'h00; mem['h2513]=8'h00;
    mem['h2514]=8'h00; mem['h2515]=8'h00; mem['h2516]=8'h00; mem['h2517]=8'h00;
    mem['h2518]=8'h00; mem['h2519]=8'h00; mem['h251A]=8'h00; mem['h251B]=8'h00;
    mem['h251C]=8'h00; mem['h251D]=8'h00; mem['h251E]=8'h00; mem['h251F]=8'h00;
    mem['h2520]=8'h00; mem['h2521]=8'h00; mem['h2522]=8'h00; mem['h2523]=8'h00;
    mem['h2524]=8'h00; mem['h2525]=8'h00; mem['h2526]=8'h00; mem['h2527]=8'h00;
    mem['h2528]=8'h00; mem['h2529]=8'h00; mem['h252A]=8'h00; mem['h252B]=8'h00;
    mem['h252C]=8'h00; mem['h252D]=8'h00; mem['h252E]=8'h00; mem['h252F]=8'h00;
    mem['h2530]=8'h00; mem['h2531]=8'h00; mem['h2532]=8'h00; mem['h2533]=8'h00;
    mem['h2534]=8'h00; mem['h2535]=8'h00; mem['h2536]=8'h00; mem['h2537]=8'h00;
    mem['h2538]=8'h00; mem['h2539]=8'h00; mem['h253A]=8'h00; mem['h253B]=8'h00;
    mem['h253C]=8'h00; mem['h253D]=8'h00; mem['h253E]=8'h00; mem['h253F]=8'h00;
    mem['h2540]=8'h00; mem['h2541]=8'h00; mem['h2542]=8'h00; mem['h2543]=8'h00;
    mem['h2544]=8'h00; mem['h2545]=8'h00; mem['h2546]=8'h00; mem['h2547]=8'h00;
    mem['h2548]=8'h00; mem['h2549]=8'h00; mem['h254A]=8'h00; mem['h254B]=8'h00;
    mem['h254C]=8'h00; mem['h254D]=8'h00; mem['h254E]=8'h00; mem['h254F]=8'h00;
    mem['h2550]=8'h00; mem['h2551]=8'h00; mem['h2552]=8'h00; mem['h2553]=8'h00;
    mem['h2554]=8'h00; mem['h2555]=8'h00; mem['h2556]=8'h00; mem['h2557]=8'h00;
    mem['h2558]=8'h00; mem['h2559]=8'h00; mem['h255A]=8'h00; mem['h255B]=8'h00;
    mem['h255C]=8'h00; mem['h255D]=8'h00; mem['h255E]=8'h00; mem['h255F]=8'h00;
    mem['h2560]=8'h00; mem['h2561]=8'h00; mem['h2562]=8'h00; mem['h2563]=8'h00;
    mem['h2564]=8'h00; mem['h2565]=8'h00; mem['h2566]=8'h00; mem['h2567]=8'h00;
    mem['h2568]=8'h00; mem['h2569]=8'h00; mem['h256A]=8'h00; mem['h256B]=8'h00;
    mem['h256C]=8'h00; mem['h256D]=8'h00; mem['h256E]=8'h00; mem['h256F]=8'h00;
    mem['h2570]=8'h00; mem['h2571]=8'h00; mem['h2572]=8'h00; mem['h2573]=8'h00;
    mem['h2574]=8'h00; mem['h2575]=8'h00; mem['h2576]=8'h00; mem['h2577]=8'h00;
    mem['h2578]=8'h00; mem['h2579]=8'h00; mem['h257A]=8'h00; mem['h257B]=8'h00;
    mem['h257C]=8'h00; mem['h257D]=8'h00; mem['h257E]=8'h00; mem['h257F]=8'h00;
    mem['h2580]=8'h00; mem['h2581]=8'h00; mem['h2582]=8'h00; mem['h2583]=8'h00;
    mem['h2584]=8'h00; mem['h2585]=8'h00; mem['h2586]=8'h00; mem['h2587]=8'h00;
    mem['h2588]=8'h00; mem['h2589]=8'h00; mem['h258A]=8'h00; mem['h258B]=8'h00;
    mem['h258C]=8'h00; mem['h258D]=8'h00; mem['h258E]=8'h00; mem['h258F]=8'h00;
    mem['h2590]=8'h00; mem['h2591]=8'h00; mem['h2592]=8'h00; mem['h2593]=8'h00;
    mem['h2594]=8'h00; mem['h2595]=8'h00; mem['h2596]=8'h00; mem['h2597]=8'h00;
    mem['h2598]=8'h00; mem['h2599]=8'h00; mem['h259A]=8'h00; mem['h259B]=8'h00;
    mem['h259C]=8'h00; mem['h259D]=8'h00; mem['h259E]=8'h00; mem['h259F]=8'h00;
    mem['h25A0]=8'h00; mem['h25A1]=8'h00; mem['h25A2]=8'h00; mem['h25A3]=8'h00;
    mem['h25A4]=8'h00; mem['h25A5]=8'h00; mem['h25A6]=8'h00; mem['h25A7]=8'h00;
    mem['h25A8]=8'h00; mem['h25A9]=8'h00; mem['h25AA]=8'h00; mem['h25AB]=8'h00;
    mem['h25AC]=8'h00; mem['h25AD]=8'h00; mem['h25AE]=8'h00; mem['h25AF]=8'h00;
    mem['h25B0]=8'h00; mem['h25B1]=8'h00; mem['h25B2]=8'h00; mem['h25B3]=8'h00;
    mem['h25B4]=8'h00; mem['h25B5]=8'h00; mem['h25B6]=8'h00; mem['h25B7]=8'h00;
    mem['h25B8]=8'h00; mem['h25B9]=8'h00; mem['h25BA]=8'h00; mem['h25BB]=8'h00;
    mem['h25BC]=8'h00; mem['h25BD]=8'h00; mem['h25BE]=8'h00; mem['h25BF]=8'h00;
    mem['h25C0]=8'h00; mem['h25C1]=8'h00; mem['h25C2]=8'h00; mem['h25C3]=8'h00;
    mem['h25C4]=8'h00; mem['h25C5]=8'h00; mem['h25C6]=8'h00; mem['h25C7]=8'h00;
    mem['h25C8]=8'h00; mem['h25C9]=8'h00; mem['h25CA]=8'h00; mem['h25CB]=8'h00;
    mem['h25CC]=8'h00; mem['h25CD]=8'h00; mem['h25CE]=8'h00; mem['h25CF]=8'h00;
    mem['h25D0]=8'h00; mem['h25D1]=8'h00; mem['h25D2]=8'h00; mem['h25D3]=8'h00;
    mem['h25D4]=8'h00; mem['h25D5]=8'h00; mem['h25D6]=8'h00; mem['h25D7]=8'h00;
    mem['h25D8]=8'h00; mem['h25D9]=8'h00; mem['h25DA]=8'h00; mem['h25DB]=8'h00;
    mem['h25DC]=8'h00; mem['h25DD]=8'h00; mem['h25DE]=8'h00; mem['h25DF]=8'h00;
    mem['h25E0]=8'h00; mem['h25E1]=8'h00; mem['h25E2]=8'h00; mem['h25E3]=8'h00;
    mem['h25E4]=8'h00; mem['h25E5]=8'h00; mem['h25E6]=8'h00; mem['h25E7]=8'h00;
    mem['h25E8]=8'h00; mem['h25E9]=8'h00; mem['h25EA]=8'h00; mem['h25EB]=8'h00;
    mem['h25EC]=8'h00; mem['h25ED]=8'h00; mem['h25EE]=8'h00; mem['h25EF]=8'h00;
    mem['h25F0]=8'h00; mem['h25F1]=8'h00; mem['h25F2]=8'h00; mem['h25F3]=8'h00;
    mem['h25F4]=8'h00; mem['h25F5]=8'h00; mem['h25F6]=8'h00; mem['h25F7]=8'h00;
    mem['h25F8]=8'h00; mem['h25F9]=8'h00; mem['h25FA]=8'h00; mem['h25FB]=8'h00;
    mem['h25FC]=8'h00; mem['h25FD]=8'h00; mem['h25FE]=8'h00; mem['h25FF]=8'h00;
    mem['h2600]=8'h00; mem['h2601]=8'h00; mem['h2602]=8'h00; mem['h2603]=8'h00;
    mem['h2604]=8'h00; mem['h2605]=8'h00; mem['h2606]=8'h00; mem['h2607]=8'h00;
    mem['h2608]=8'h00; mem['h2609]=8'h00; mem['h260A]=8'h00; mem['h260B]=8'h00;
    mem['h260C]=8'h00; mem['h260D]=8'h00; mem['h260E]=8'h00; mem['h260F]=8'h00;
    mem['h2610]=8'h00; mem['h2611]=8'h00; mem['h2612]=8'h00; mem['h2613]=8'h00;
    mem['h2614]=8'h00; mem['h2615]=8'h00; mem['h2616]=8'h00; mem['h2617]=8'h00;
    mem['h2618]=8'h00; mem['h2619]=8'h00; mem['h261A]=8'h00; mem['h261B]=8'h00;
    mem['h261C]=8'h00; mem['h261D]=8'h00; mem['h261E]=8'h00; mem['h261F]=8'h00;
    mem['h2620]=8'h00; mem['h2621]=8'h00; mem['h2622]=8'h00; mem['h2623]=8'h00;
    mem['h2624]=8'h00; mem['h2625]=8'h00; mem['h2626]=8'h00; mem['h2627]=8'h00;
    mem['h2628]=8'h00; mem['h2629]=8'h00; mem['h262A]=8'h00; mem['h262B]=8'h00;
    mem['h262C]=8'h00; mem['h262D]=8'h00; mem['h262E]=8'h00; mem['h262F]=8'h00;
    mem['h2630]=8'h00; mem['h2631]=8'h00; mem['h2632]=8'h00; mem['h2633]=8'h00;
    mem['h2634]=8'h00; mem['h2635]=8'h00; mem['h2636]=8'h00; mem['h2637]=8'h00;
    mem['h2638]=8'h00; mem['h2639]=8'h00; mem['h263A]=8'h00; mem['h263B]=8'h00;
    mem['h263C]=8'h00; mem['h263D]=8'h00; mem['h263E]=8'h00; mem['h263F]=8'h00;
    mem['h2640]=8'h00; mem['h2641]=8'h00; mem['h2642]=8'h00; mem['h2643]=8'h00;
    mem['h2644]=8'h00; mem['h2645]=8'h00; mem['h2646]=8'h00; mem['h2647]=8'h00;
    mem['h2648]=8'h00; mem['h2649]=8'h00; mem['h264A]=8'h00; mem['h264B]=8'h00;
    mem['h264C]=8'h00; mem['h264D]=8'h00; mem['h264E]=8'h00; mem['h264F]=8'h00;
    mem['h2650]=8'h00; mem['h2651]=8'h00; mem['h2652]=8'h00; mem['h2653]=8'h00;
    mem['h2654]=8'h00; mem['h2655]=8'h00; mem['h2656]=8'h00; mem['h2657]=8'h00;
    mem['h2658]=8'h00; mem['h2659]=8'h00; mem['h265A]=8'h00; mem['h265B]=8'h00;
    mem['h265C]=8'h00; mem['h265D]=8'h00; mem['h265E]=8'h00; mem['h265F]=8'h00;
    mem['h2660]=8'h00; mem['h2661]=8'h00; mem['h2662]=8'h00; mem['h2663]=8'h00;
    mem['h2664]=8'h00; mem['h2665]=8'h00; mem['h2666]=8'h00; mem['h2667]=8'h00;
    mem['h2668]=8'h00; mem['h2669]=8'h00; mem['h266A]=8'h00; mem['h266B]=8'h00;
    mem['h266C]=8'h00; mem['h266D]=8'h00; mem['h266E]=8'h00; mem['h266F]=8'h00;
    mem['h2670]=8'h00; mem['h2671]=8'h00; mem['h2672]=8'h00; mem['h2673]=8'h00;
    mem['h2674]=8'h00; mem['h2675]=8'h00; mem['h2676]=8'h00; mem['h2677]=8'h00;
    mem['h2678]=8'h00; mem['h2679]=8'h00; mem['h267A]=8'h00; mem['h267B]=8'h00;
    mem['h267C]=8'h00; mem['h267D]=8'h00; mem['h267E]=8'h00; mem['h267F]=8'h00;
    mem['h2680]=8'h00; mem['h2681]=8'h00; mem['h2682]=8'h00; mem['h2683]=8'h00;
    mem['h2684]=8'h00; mem['h2685]=8'h00; mem['h2686]=8'h00; mem['h2687]=8'h00;
    mem['h2688]=8'h00; mem['h2689]=8'h00; mem['h268A]=8'h00; mem['h268B]=8'h00;
    mem['h268C]=8'h00; mem['h268D]=8'h00; mem['h268E]=8'h00; mem['h268F]=8'h00;
    mem['h2690]=8'h00; mem['h2691]=8'h00; mem['h2692]=8'h00; mem['h2693]=8'h00;
    mem['h2694]=8'h00; mem['h2695]=8'h00; mem['h2696]=8'h00; mem['h2697]=8'h00;
    mem['h2698]=8'h00; mem['h2699]=8'h00; mem['h269A]=8'h00; mem['h269B]=8'h00;
    mem['h269C]=8'h00; mem['h269D]=8'h00; mem['h269E]=8'h00; mem['h269F]=8'h00;
    mem['h26A0]=8'h00; mem['h26A1]=8'h00; mem['h26A2]=8'h00; mem['h26A3]=8'h00;
    mem['h26A4]=8'h00; mem['h26A5]=8'h00; mem['h26A6]=8'h00; mem['h26A7]=8'h00;
    mem['h26A8]=8'h00; mem['h26A9]=8'h00; mem['h26AA]=8'h00; mem['h26AB]=8'h00;
    mem['h26AC]=8'h00; mem['h26AD]=8'h00; mem['h26AE]=8'h00; mem['h26AF]=8'h00;
    mem['h26B0]=8'h00; mem['h26B1]=8'h00; mem['h26B2]=8'h00; mem['h26B3]=8'h00;
    mem['h26B4]=8'h00; mem['h26B5]=8'h00; mem['h26B6]=8'h00; mem['h26B7]=8'h00;
    mem['h26B8]=8'h00; mem['h26B9]=8'h00; mem['h26BA]=8'h00; mem['h26BB]=8'h00;
    mem['h26BC]=8'h00; mem['h26BD]=8'h00; mem['h26BE]=8'h00; mem['h26BF]=8'h00;
    mem['h26C0]=8'h00; mem['h26C1]=8'h00; mem['h26C2]=8'h00; mem['h26C3]=8'h00;
    mem['h26C4]=8'h00; mem['h26C5]=8'h00; mem['h26C6]=8'h00; mem['h26C7]=8'h00;
    mem['h26C8]=8'h00; mem['h26C9]=8'h00; mem['h26CA]=8'h00; mem['h26CB]=8'h00;
    mem['h26CC]=8'h00; mem['h26CD]=8'h00; mem['h26CE]=8'h00; mem['h26CF]=8'h00;
    mem['h26D0]=8'h00; mem['h26D1]=8'h00; mem['h26D2]=8'h00; mem['h26D3]=8'h00;
    mem['h26D4]=8'h00; mem['h26D5]=8'h00; mem['h26D6]=8'h00; mem['h26D7]=8'h00;
    mem['h26D8]=8'h00; mem['h26D9]=8'h00; mem['h26DA]=8'h00; mem['h26DB]=8'h00;
    mem['h26DC]=8'h00; mem['h26DD]=8'h00; mem['h26DE]=8'h00; mem['h26DF]=8'h00;
    mem['h26E0]=8'h00; mem['h26E1]=8'h00; mem['h26E2]=8'h00; mem['h26E3]=8'h00;
    mem['h26E4]=8'h00; mem['h26E5]=8'h00; mem['h26E6]=8'h00; mem['h26E7]=8'h00;
    mem['h26E8]=8'h00; mem['h26E9]=8'h00; mem['h26EA]=8'h00; mem['h26EB]=8'h00;
    mem['h26EC]=8'h00; mem['h26ED]=8'h00; mem['h26EE]=8'h00; mem['h26EF]=8'h00;
    mem['h26F0]=8'h00; mem['h26F1]=8'h00; mem['h26F2]=8'h00; mem['h26F3]=8'h00;
    mem['h26F4]=8'h00; mem['h26F5]=8'h00; mem['h26F6]=8'h00; mem['h26F7]=8'h00;
    mem['h26F8]=8'h00; mem['h26F9]=8'h00; mem['h26FA]=8'h00; mem['h26FB]=8'h00;
    mem['h26FC]=8'h00; mem['h26FD]=8'h00; mem['h26FE]=8'h00; mem['h26FF]=8'h00;
    mem['h2700]=8'h00; mem['h2701]=8'h00; mem['h2702]=8'h00; mem['h2703]=8'h00;
    mem['h2704]=8'h00; mem['h2705]=8'h00; mem['h2706]=8'h00; mem['h2707]=8'h00;
    mem['h2708]=8'h00; mem['h2709]=8'h00; mem['h270A]=8'h00; mem['h270B]=8'h00;
    mem['h270C]=8'h00; mem['h270D]=8'h00; mem['h270E]=8'h00; mem['h270F]=8'h00;
    mem['h2710]=8'h00; mem['h2711]=8'h00; mem['h2712]=8'h00; mem['h2713]=8'h00;
    mem['h2714]=8'h00; mem['h2715]=8'h00; mem['h2716]=8'h00; mem['h2717]=8'h00;
    mem['h2718]=8'h00; mem['h2719]=8'h00; mem['h271A]=8'h00; mem['h271B]=8'h00;
    mem['h271C]=8'h00; mem['h271D]=8'h00; mem['h271E]=8'h00; mem['h271F]=8'h00;
    mem['h2720]=8'h00; mem['h2721]=8'h00; mem['h2722]=8'h00; mem['h2723]=8'h00;
    mem['h2724]=8'h00; mem['h2725]=8'h00; mem['h2726]=8'h00; mem['h2727]=8'h00;
    mem['h2728]=8'h00; mem['h2729]=8'h00; mem['h272A]=8'h00; mem['h272B]=8'h00;
    mem['h272C]=8'h00; mem['h272D]=8'h00; mem['h272E]=8'h00; mem['h272F]=8'h00;
    mem['h2730]=8'h00; mem['h2731]=8'h00; mem['h2732]=8'h00; mem['h2733]=8'h00;
    mem['h2734]=8'h00; mem['h2735]=8'h00; mem['h2736]=8'h00; mem['h2737]=8'h00;
    mem['h2738]=8'h00; mem['h2739]=8'h00; mem['h273A]=8'h00; mem['h273B]=8'h00;
    mem['h273C]=8'h00; mem['h273D]=8'h00; mem['h273E]=8'h00; mem['h273F]=8'h00;
    mem['h2740]=8'h00; mem['h2741]=8'h00; mem['h2742]=8'h00; mem['h2743]=8'h00;
    mem['h2744]=8'h00; mem['h2745]=8'h00; mem['h2746]=8'h00; mem['h2747]=8'h00;
    mem['h2748]=8'h00; mem['h2749]=8'h00; mem['h274A]=8'h00; mem['h274B]=8'h00;
    mem['h274C]=8'h00; mem['h274D]=8'h00; mem['h274E]=8'h00; mem['h274F]=8'h00;
    mem['h2750]=8'h00; mem['h2751]=8'h00; mem['h2752]=8'h00; mem['h2753]=8'h00;
    mem['h2754]=8'h00; mem['h2755]=8'h00; mem['h2756]=8'h00; mem['h2757]=8'h00;
    mem['h2758]=8'h00; mem['h2759]=8'h00; mem['h275A]=8'h00; mem['h275B]=8'h00;
    mem['h275C]=8'h00; mem['h275D]=8'h00; mem['h275E]=8'h00; mem['h275F]=8'h00;
    mem['h2760]=8'h00; mem['h2761]=8'h00; mem['h2762]=8'h00; mem['h2763]=8'h00;
    mem['h2764]=8'h00; mem['h2765]=8'h00; mem['h2766]=8'h00; mem['h2767]=8'h00;
    mem['h2768]=8'h00; mem['h2769]=8'h00; mem['h276A]=8'h00; mem['h276B]=8'h00;
    mem['h276C]=8'h00; mem['h276D]=8'h00; mem['h276E]=8'h00; mem['h276F]=8'h00;
    mem['h2770]=8'h00; mem['h2771]=8'h00; mem['h2772]=8'h00; mem['h2773]=8'h00;
    mem['h2774]=8'h00; mem['h2775]=8'h00; mem['h2776]=8'h00; mem['h2777]=8'h00;
    mem['h2778]=8'h00; mem['h2779]=8'h00; mem['h277A]=8'h00; mem['h277B]=8'h00;
    mem['h277C]=8'h00; mem['h277D]=8'h00; mem['h277E]=8'h00; mem['h277F]=8'h00;
    mem['h2780]=8'h00; mem['h2781]=8'h00; mem['h2782]=8'h00; mem['h2783]=8'h00;
    mem['h2784]=8'h00; mem['h2785]=8'h00; mem['h2786]=8'h00; mem['h2787]=8'h00;
    mem['h2788]=8'h00; mem['h2789]=8'h00; mem['h278A]=8'h00; mem['h278B]=8'h00;
    mem['h278C]=8'h00; mem['h278D]=8'h00; mem['h278E]=8'h00; mem['h278F]=8'h00;
    mem['h2790]=8'h00; mem['h2791]=8'h00; mem['h2792]=8'h00; mem['h2793]=8'h00;
    mem['h2794]=8'h00; mem['h2795]=8'h00; mem['h2796]=8'h00; mem['h2797]=8'h00;
    mem['h2798]=8'h00; mem['h2799]=8'h00; mem['h279A]=8'h00; mem['h279B]=8'h00;
    mem['h279C]=8'h00; mem['h279D]=8'h00; mem['h279E]=8'h00; mem['h279F]=8'h00;
    mem['h27A0]=8'h00; mem['h27A1]=8'h00; mem['h27A2]=8'h00; mem['h27A3]=8'h00;
    mem['h27A4]=8'h00; mem['h27A5]=8'h00; mem['h27A6]=8'h00; mem['h27A7]=8'h00;
    mem['h27A8]=8'h00; mem['h27A9]=8'h00; mem['h27AA]=8'h00; mem['h27AB]=8'h00;
    mem['h27AC]=8'h00; mem['h27AD]=8'h00; mem['h27AE]=8'h00; mem['h27AF]=8'h00;
    mem['h27B0]=8'h00; mem['h27B1]=8'h00; mem['h27B2]=8'h00; mem['h27B3]=8'h00;
    mem['h27B4]=8'h00; mem['h27B5]=8'h00; mem['h27B6]=8'h00; mem['h27B7]=8'h00;
    mem['h27B8]=8'h00; mem['h27B9]=8'h00; mem['h27BA]=8'h00; mem['h27BB]=8'h00;
    mem['h27BC]=8'h00; mem['h27BD]=8'h00; mem['h27BE]=8'h00; mem['h27BF]=8'h00;
    mem['h27C0]=8'h00; mem['h27C1]=8'h00; mem['h27C2]=8'h00; mem['h27C3]=8'h00;
    mem['h27C4]=8'h00; mem['h27C5]=8'h00; mem['h27C6]=8'h00; mem['h27C7]=8'h00;
    mem['h27C8]=8'h00; mem['h27C9]=8'h00; mem['h27CA]=8'h00; mem['h27CB]=8'h00;
    mem['h27CC]=8'h00; mem['h27CD]=8'h00; mem['h27CE]=8'h00; mem['h27CF]=8'h00;
    mem['h27D0]=8'h00; mem['h27D1]=8'h00; mem['h27D2]=8'h00; mem['h27D3]=8'h00;
    mem['h27D4]=8'h00; mem['h27D5]=8'h00; mem['h27D6]=8'h00; mem['h27D7]=8'h00;
    mem['h27D8]=8'h00; mem['h27D9]=8'h00; mem['h27DA]=8'h00; mem['h27DB]=8'h00;
    mem['h27DC]=8'h00; mem['h27DD]=8'h00; mem['h27DE]=8'h00; mem['h27DF]=8'h00;
    mem['h27E0]=8'h00; mem['h27E1]=8'h00; mem['h27E2]=8'h00; mem['h27E3]=8'h00;
    mem['h27E4]=8'h00; mem['h27E5]=8'h00; mem['h27E6]=8'h00; mem['h27E7]=8'h00;
    mem['h27E8]=8'h00; mem['h27E9]=8'h00; mem['h27EA]=8'h00; mem['h27EB]=8'h00;
    mem['h27EC]=8'h00; mem['h27ED]=8'h00; mem['h27EE]=8'h00; mem['h27EF]=8'h00;
    mem['h27F0]=8'h00; mem['h27F1]=8'h00; mem['h27F2]=8'h00; mem['h27F3]=8'h00;
    mem['h27F4]=8'h00; mem['h27F5]=8'h00; mem['h27F6]=8'h00; mem['h27F7]=8'h00;
    mem['h27F8]=8'h00; mem['h27F9]=8'h00; mem['h27FA]=8'h00; mem['h27FB]=8'h00;
    mem['h27FC]=8'h00; mem['h27FD]=8'h00; mem['h27FE]=8'h00; mem['h27FF]=8'h00;
    mem['h2800]=8'h00; mem['h2801]=8'h00; mem['h2802]=8'h00; mem['h2803]=8'h00;
    mem['h2804]=8'h00; mem['h2805]=8'h00; mem['h2806]=8'h00; mem['h2807]=8'h00;
    mem['h2808]=8'h00; mem['h2809]=8'h00; mem['h280A]=8'h00; mem['h280B]=8'h00;
    mem['h280C]=8'h00; mem['h280D]=8'h00; mem['h280E]=8'h00; mem['h280F]=8'h00;
    mem['h2810]=8'h00; mem['h2811]=8'h00; mem['h2812]=8'h00; mem['h2813]=8'h00;
    mem['h2814]=8'h00; mem['h2815]=8'h00; mem['h2816]=8'h00; mem['h2817]=8'h00;
    mem['h2818]=8'h00; mem['h2819]=8'h00; mem['h281A]=8'h00; mem['h281B]=8'h00;
    mem['h281C]=8'h00; mem['h281D]=8'h00; mem['h281E]=8'h00; mem['h281F]=8'h00;
    mem['h2820]=8'h00; mem['h2821]=8'h00; mem['h2822]=8'h00; mem['h2823]=8'h00;
    mem['h2824]=8'h00; mem['h2825]=8'h00; mem['h2826]=8'h00; mem['h2827]=8'h00;
    mem['h2828]=8'h00; mem['h2829]=8'h00; mem['h282A]=8'h00; mem['h282B]=8'h00;
    mem['h282C]=8'h00; mem['h282D]=8'h00; mem['h282E]=8'h00; mem['h282F]=8'h00;
    mem['h2830]=8'h00; mem['h2831]=8'h00; mem['h2832]=8'h00; mem['h2833]=8'h00;
    mem['h2834]=8'h00; mem['h2835]=8'h00; mem['h2836]=8'h00; mem['h2837]=8'h00;
    mem['h2838]=8'h00; mem['h2839]=8'h00; mem['h283A]=8'h00; mem['h283B]=8'h00;
    mem['h283C]=8'h00; mem['h283D]=8'h00; mem['h283E]=8'h00; mem['h283F]=8'h00;
    mem['h2840]=8'h00; mem['h2841]=8'h00; mem['h2842]=8'h00; mem['h2843]=8'h00;
    mem['h2844]=8'h00; mem['h2845]=8'h00; mem['h2846]=8'h00; mem['h2847]=8'h00;
    mem['h2848]=8'h00; mem['h2849]=8'h00; mem['h284A]=8'h00; mem['h284B]=8'h00;
    mem['h284C]=8'h00; mem['h284D]=8'h00; mem['h284E]=8'h00; mem['h284F]=8'h00;
    mem['h2850]=8'h00; mem['h2851]=8'h00; mem['h2852]=8'h00; mem['h2853]=8'h00;
    mem['h2854]=8'h00; mem['h2855]=8'h00; mem['h2856]=8'h00; mem['h2857]=8'h00;
    mem['h2858]=8'h00; mem['h2859]=8'h00; mem['h285A]=8'h00; mem['h285B]=8'h00;
    mem['h285C]=8'h00; mem['h285D]=8'h00; mem['h285E]=8'h00; mem['h285F]=8'h00;
    mem['h2860]=8'h00; mem['h2861]=8'h00; mem['h2862]=8'h00; mem['h2863]=8'h00;
    mem['h2864]=8'h00; mem['h2865]=8'h00; mem['h2866]=8'h00; mem['h2867]=8'h00;
    mem['h2868]=8'h00; mem['h2869]=8'h00; mem['h286A]=8'h00; mem['h286B]=8'h00;
    mem['h286C]=8'h00; mem['h286D]=8'h00; mem['h286E]=8'h00; mem['h286F]=8'h00;
    mem['h2870]=8'h00; mem['h2871]=8'h00; mem['h2872]=8'h00; mem['h2873]=8'h00;
    mem['h2874]=8'h00; mem['h2875]=8'h00; mem['h2876]=8'h00; mem['h2877]=8'h00;
    mem['h2878]=8'h00; mem['h2879]=8'h00; mem['h287A]=8'h00; mem['h287B]=8'h00;
    mem['h287C]=8'h00; mem['h287D]=8'h00; mem['h287E]=8'h00; mem['h287F]=8'h00;
    mem['h2880]=8'h00; mem['h2881]=8'h00; mem['h2882]=8'h00; mem['h2883]=8'h00;
    mem['h2884]=8'h00; mem['h2885]=8'h00; mem['h2886]=8'h00; mem['h2887]=8'h00;
    mem['h2888]=8'h00; mem['h2889]=8'h00; mem['h288A]=8'h00; mem['h288B]=8'h00;
    mem['h288C]=8'h00; mem['h288D]=8'h00; mem['h288E]=8'h00; mem['h288F]=8'h00;
    mem['h2890]=8'h00; mem['h2891]=8'h00; mem['h2892]=8'h00; mem['h2893]=8'h00;
    mem['h2894]=8'h00; mem['h2895]=8'h00; mem['h2896]=8'h00; mem['h2897]=8'h00;
    mem['h2898]=8'h00; mem['h2899]=8'h00; mem['h289A]=8'h00; mem['h289B]=8'h00;
    mem['h289C]=8'h00; mem['h289D]=8'h00; mem['h289E]=8'h00; mem['h289F]=8'h00;
    mem['h28A0]=8'h00; mem['h28A1]=8'h00; mem['h28A2]=8'h00; mem['h28A3]=8'h00;
    mem['h28A4]=8'h00; mem['h28A5]=8'h00; mem['h28A6]=8'h00; mem['h28A7]=8'h00;
    mem['h28A8]=8'h00; mem['h28A9]=8'h00; mem['h28AA]=8'h00; mem['h28AB]=8'h00;
    mem['h28AC]=8'h00; mem['h28AD]=8'h00; mem['h28AE]=8'h00; mem['h28AF]=8'h00;
    mem['h28B0]=8'h00; mem['h28B1]=8'h00; mem['h28B2]=8'h00; mem['h28B3]=8'h00;
    mem['h28B4]=8'h00; mem['h28B5]=8'h00; mem['h28B6]=8'h00; mem['h28B7]=8'h00;
    mem['h28B8]=8'h00; mem['h28B9]=8'h00; mem['h28BA]=8'h00; mem['h28BB]=8'h00;
    mem['h28BC]=8'h00; mem['h28BD]=8'h00; mem['h28BE]=8'h00; mem['h28BF]=8'h00;
    mem['h28C0]=8'h00; mem['h28C1]=8'h00; mem['h28C2]=8'h00; mem['h28C3]=8'h00;
    mem['h28C4]=8'h00; mem['h28C5]=8'h00; mem['h28C6]=8'h00; mem['h28C7]=8'h00;
    mem['h28C8]=8'h00; mem['h28C9]=8'h00; mem['h28CA]=8'h00; mem['h28CB]=8'h00;
    mem['h28CC]=8'h00; mem['h28CD]=8'h00; mem['h28CE]=8'h00; mem['h28CF]=8'h00;
    mem['h28D0]=8'h00; mem['h28D1]=8'h00; mem['h28D2]=8'h00; mem['h28D3]=8'h00;
    mem['h28D4]=8'h00; mem['h28D5]=8'h00; mem['h28D6]=8'h00; mem['h28D7]=8'h00;
    mem['h28D8]=8'h00; mem['h28D9]=8'h00; mem['h28DA]=8'h00; mem['h28DB]=8'h00;
    mem['h28DC]=8'h00; mem['h28DD]=8'h00; mem['h28DE]=8'h00; mem['h28DF]=8'h00;
    mem['h28E0]=8'h00; mem['h28E1]=8'h00; mem['h28E2]=8'h00; mem['h28E3]=8'h00;
    mem['h28E4]=8'h00; mem['h28E5]=8'h00; mem['h28E6]=8'h00; mem['h28E7]=8'h00;
    mem['h28E8]=8'h00; mem['h28E9]=8'h00; mem['h28EA]=8'h00; mem['h28EB]=8'h00;
    mem['h28EC]=8'h00; mem['h28ED]=8'h00; mem['h28EE]=8'h00; mem['h28EF]=8'h00;
    mem['h28F0]=8'h00; mem['h28F1]=8'h00; mem['h28F2]=8'h00; mem['h28F3]=8'h00;
    mem['h28F4]=8'h00; mem['h28F5]=8'h00; mem['h28F6]=8'h00; mem['h28F7]=8'h00;
    mem['h28F8]=8'h00; mem['h28F9]=8'h00; mem['h28FA]=8'h00; mem['h28FB]=8'h00;
    mem['h28FC]=8'h00; mem['h28FD]=8'h00; mem['h28FE]=8'h00; mem['h28FF]=8'h00;
    mem['h2900]=8'h00; mem['h2901]=8'h00; mem['h2902]=8'h00; mem['h2903]=8'h00;
    mem['h2904]=8'h00; mem['h2905]=8'h00; mem['h2906]=8'h00; mem['h2907]=8'h00;
    mem['h2908]=8'h00; mem['h2909]=8'h00; mem['h290A]=8'h00; mem['h290B]=8'h00;
    mem['h290C]=8'h00; mem['h290D]=8'h00; mem['h290E]=8'h00; mem['h290F]=8'h00;
    mem['h2910]=8'h00; mem['h2911]=8'h00; mem['h2912]=8'h00; mem['h2913]=8'h00;
    mem['h2914]=8'h00; mem['h2915]=8'h00; mem['h2916]=8'h00; mem['h2917]=8'h00;
    mem['h2918]=8'h00; mem['h2919]=8'h00; mem['h291A]=8'h00; mem['h291B]=8'h00;
    mem['h291C]=8'h00; mem['h291D]=8'h00; mem['h291E]=8'h00; mem['h291F]=8'h00;
    mem['h2920]=8'h00; mem['h2921]=8'h00; mem['h2922]=8'h00; mem['h2923]=8'h00;
    mem['h2924]=8'h00; mem['h2925]=8'h00; mem['h2926]=8'h00; mem['h2927]=8'h00;
    mem['h2928]=8'h00; mem['h2929]=8'h00; mem['h292A]=8'h00; mem['h292B]=8'h00;
    mem['h292C]=8'h00; mem['h292D]=8'h00; mem['h292E]=8'h00; mem['h292F]=8'h00;
    mem['h2930]=8'h00; mem['h2931]=8'h00; mem['h2932]=8'h00; mem['h2933]=8'h00;
    mem['h2934]=8'h00; mem['h2935]=8'h00; mem['h2936]=8'h00; mem['h2937]=8'h00;
    mem['h2938]=8'h00; mem['h2939]=8'h00; mem['h293A]=8'h00; mem['h293B]=8'h00;
    mem['h293C]=8'h00; mem['h293D]=8'h00; mem['h293E]=8'h00; mem['h293F]=8'h00;
    mem['h2940]=8'h00; mem['h2941]=8'h00; mem['h2942]=8'h00; mem['h2943]=8'h00;
    mem['h2944]=8'h00; mem['h2945]=8'h00; mem['h2946]=8'h00; mem['h2947]=8'h00;
    mem['h2948]=8'h00; mem['h2949]=8'h00; mem['h294A]=8'h00; mem['h294B]=8'h00;
    mem['h294C]=8'h00; mem['h294D]=8'h00; mem['h294E]=8'h00; mem['h294F]=8'h00;
    mem['h2950]=8'h00; mem['h2951]=8'h00; mem['h2952]=8'h00; mem['h2953]=8'h00;
    mem['h2954]=8'h00; mem['h2955]=8'h00; mem['h2956]=8'h00; mem['h2957]=8'h00;
    mem['h2958]=8'h00; mem['h2959]=8'h00; mem['h295A]=8'h00; mem['h295B]=8'h00;
    mem['h295C]=8'h00; mem['h295D]=8'h00; mem['h295E]=8'h00; mem['h295F]=8'h00;
    mem['h2960]=8'h00; mem['h2961]=8'h00; mem['h2962]=8'h00; mem['h2963]=8'h00;
    mem['h2964]=8'h00; mem['h2965]=8'h00; mem['h2966]=8'h00; mem['h2967]=8'h00;
    mem['h2968]=8'h00; mem['h2969]=8'h00; mem['h296A]=8'h00; mem['h296B]=8'h00;
    mem['h296C]=8'h00; mem['h296D]=8'h00; mem['h296E]=8'h00; mem['h296F]=8'h00;
    mem['h2970]=8'h00; mem['h2971]=8'h00; mem['h2972]=8'h00; mem['h2973]=8'h00;
    mem['h2974]=8'h00; mem['h2975]=8'h00; mem['h2976]=8'h00; mem['h2977]=8'h00;
    mem['h2978]=8'h00; mem['h2979]=8'h00; mem['h297A]=8'h00; mem['h297B]=8'h00;
    mem['h297C]=8'h00; mem['h297D]=8'h00; mem['h297E]=8'h00; mem['h297F]=8'h00;
    mem['h2980]=8'h00; mem['h2981]=8'h00; mem['h2982]=8'h00; mem['h2983]=8'h00;
    mem['h2984]=8'h00; mem['h2985]=8'h00; mem['h2986]=8'h00; mem['h2987]=8'h00;
    mem['h2988]=8'h00; mem['h2989]=8'h00; mem['h298A]=8'h00; mem['h298B]=8'h00;
    mem['h298C]=8'h00; mem['h298D]=8'h00; mem['h298E]=8'h00; mem['h298F]=8'h00;
    mem['h2990]=8'h00; mem['h2991]=8'h00; mem['h2992]=8'h00; mem['h2993]=8'h00;
    mem['h2994]=8'h00; mem['h2995]=8'h00; mem['h2996]=8'h00; mem['h2997]=8'h00;
    mem['h2998]=8'h00; mem['h2999]=8'h00; mem['h299A]=8'h00; mem['h299B]=8'h00;
    mem['h299C]=8'h00; mem['h299D]=8'h00; mem['h299E]=8'h00; mem['h299F]=8'h00;
    mem['h29A0]=8'h00; mem['h29A1]=8'h00; mem['h29A2]=8'h00; mem['h29A3]=8'h00;
    mem['h29A4]=8'h00; mem['h29A5]=8'h00; mem['h29A6]=8'h00; mem['h29A7]=8'h00;
    mem['h29A8]=8'h00; mem['h29A9]=8'h00; mem['h29AA]=8'h00; mem['h29AB]=8'h00;
    mem['h29AC]=8'h00; mem['h29AD]=8'h00; mem['h29AE]=8'h00; mem['h29AF]=8'h00;
    mem['h29B0]=8'h00; mem['h29B1]=8'h00; mem['h29B2]=8'h00; mem['h29B3]=8'h00;
    mem['h29B4]=8'h00; mem['h29B5]=8'h00; mem['h29B6]=8'h00; mem['h29B7]=8'h00;
    mem['h29B8]=8'h00; mem['h29B9]=8'h00; mem['h29BA]=8'h00; mem['h29BB]=8'h00;
    mem['h29BC]=8'h00; mem['h29BD]=8'h00; mem['h29BE]=8'h00; mem['h29BF]=8'h00;
    mem['h29C0]=8'h00; mem['h29C1]=8'h00; mem['h29C2]=8'h00; mem['h29C3]=8'h00;
    mem['h29C4]=8'h00; mem['h29C5]=8'h00; mem['h29C6]=8'h00; mem['h29C7]=8'h00;
    mem['h29C8]=8'h00; mem['h29C9]=8'h00; mem['h29CA]=8'h00; mem['h29CB]=8'h00;
    mem['h29CC]=8'h00; mem['h29CD]=8'h00; mem['h29CE]=8'h00; mem['h29CF]=8'h00;
    mem['h29D0]=8'h00; mem['h29D1]=8'h00; mem['h29D2]=8'h00; mem['h29D3]=8'h00;
    mem['h29D4]=8'h00; mem['h29D5]=8'h00; mem['h29D6]=8'h00; mem['h29D7]=8'h00;
    mem['h29D8]=8'h00; mem['h29D9]=8'h00; mem['h29DA]=8'h00; mem['h29DB]=8'h00;
    mem['h29DC]=8'h00; mem['h29DD]=8'h00; mem['h29DE]=8'h00; mem['h29DF]=8'h00;
    mem['h29E0]=8'h00; mem['h29E1]=8'h00; mem['h29E2]=8'h00; mem['h29E3]=8'h00;
    mem['h29E4]=8'h00; mem['h29E5]=8'h00; mem['h29E6]=8'h00; mem['h29E7]=8'h00;
    mem['h29E8]=8'h00; mem['h29E9]=8'h00; mem['h29EA]=8'h00; mem['h29EB]=8'h00;
    mem['h29EC]=8'h00; mem['h29ED]=8'h00; mem['h29EE]=8'h00; mem['h29EF]=8'h00;
    mem['h29F0]=8'h00; mem['h29F1]=8'h00; mem['h29F2]=8'h00; mem['h29F3]=8'h00;
    mem['h29F4]=8'h00; mem['h29F5]=8'h00; mem['h29F6]=8'h00; mem['h29F7]=8'h00;
    mem['h29F8]=8'h00; mem['h29F9]=8'h00; mem['h29FA]=8'h00; mem['h29FB]=8'h00;
    mem['h29FC]=8'h00; mem['h29FD]=8'h00; mem['h29FE]=8'h00; mem['h29FF]=8'h00;
    mem['h2A00]=8'h00; mem['h2A01]=8'h00; mem['h2A02]=8'h00; mem['h2A03]=8'h00;
    mem['h2A04]=8'h00; mem['h2A05]=8'h00; mem['h2A06]=8'h00; mem['h2A07]=8'h00;
    mem['h2A08]=8'h00; mem['h2A09]=8'h00; mem['h2A0A]=8'h00; mem['h2A0B]=8'h00;
    mem['h2A0C]=8'h00; mem['h2A0D]=8'h00; mem['h2A0E]=8'h00; mem['h2A0F]=8'h00;
    mem['h2A10]=8'h00; mem['h2A11]=8'h00; mem['h2A12]=8'h00; mem['h2A13]=8'h00;
    mem['h2A14]=8'h00; mem['h2A15]=8'h00; mem['h2A16]=8'h00; mem['h2A17]=8'h00;
    mem['h2A18]=8'h00; mem['h2A19]=8'h00; mem['h2A1A]=8'h00; mem['h2A1B]=8'h00;
    mem['h2A1C]=8'h00; mem['h2A1D]=8'h00; mem['h2A1E]=8'h00; mem['h2A1F]=8'h00;
    mem['h2A20]=8'h00; mem['h2A21]=8'h00; mem['h2A22]=8'h00; mem['h2A23]=8'h00;
    mem['h2A24]=8'h00; mem['h2A25]=8'h00; mem['h2A26]=8'h00; mem['h2A27]=8'h00;
    mem['h2A28]=8'h00; mem['h2A29]=8'h00; mem['h2A2A]=8'h00; mem['h2A2B]=8'h00;
    mem['h2A2C]=8'h00; mem['h2A2D]=8'h00; mem['h2A2E]=8'h00; mem['h2A2F]=8'h00;
    mem['h2A30]=8'h00; mem['h2A31]=8'h00; mem['h2A32]=8'h00; mem['h2A33]=8'h00;
    mem['h2A34]=8'h00; mem['h2A35]=8'h00; mem['h2A36]=8'h00; mem['h2A37]=8'h00;
    mem['h2A38]=8'h00; mem['h2A39]=8'h00; mem['h2A3A]=8'h00; mem['h2A3B]=8'h00;
    mem['h2A3C]=8'h00; mem['h2A3D]=8'h00; mem['h2A3E]=8'h00; mem['h2A3F]=8'h00;
    mem['h2A40]=8'h00; mem['h2A41]=8'h00; mem['h2A42]=8'h00; mem['h2A43]=8'h00;
    mem['h2A44]=8'h00; mem['h2A45]=8'h00; mem['h2A46]=8'h00; mem['h2A47]=8'h00;
    mem['h2A48]=8'h00; mem['h2A49]=8'h00; mem['h2A4A]=8'h00; mem['h2A4B]=8'h00;
    mem['h2A4C]=8'h00; mem['h2A4D]=8'h00; mem['h2A4E]=8'h00; mem['h2A4F]=8'h00;
    mem['h2A50]=8'h00; mem['h2A51]=8'h00; mem['h2A52]=8'h00; mem['h2A53]=8'h00;
    mem['h2A54]=8'h00; mem['h2A55]=8'h00; mem['h2A56]=8'h00; mem['h2A57]=8'h00;
    mem['h2A58]=8'h00; mem['h2A59]=8'h00; mem['h2A5A]=8'h00; mem['h2A5B]=8'h00;
    mem['h2A5C]=8'h00; mem['h2A5D]=8'h00; mem['h2A5E]=8'h00; mem['h2A5F]=8'h00;
    mem['h2A60]=8'h00; mem['h2A61]=8'h00; mem['h2A62]=8'h00; mem['h2A63]=8'h00;
    mem['h2A64]=8'h00; mem['h2A65]=8'h00; mem['h2A66]=8'h00; mem['h2A67]=8'h00;
    mem['h2A68]=8'h00; mem['h2A69]=8'h00; mem['h2A6A]=8'h00; mem['h2A6B]=8'h00;
    mem['h2A6C]=8'h00; mem['h2A6D]=8'h00; mem['h2A6E]=8'h00; mem['h2A6F]=8'h00;
    mem['h2A70]=8'h00; mem['h2A71]=8'h00; mem['h2A72]=8'h00; mem['h2A73]=8'h00;
    mem['h2A74]=8'h00; mem['h2A75]=8'h00; mem['h2A76]=8'h00; mem['h2A77]=8'h00;
    mem['h2A78]=8'h00; mem['h2A79]=8'h00; mem['h2A7A]=8'h00; mem['h2A7B]=8'h00;
    mem['h2A7C]=8'h00; mem['h2A7D]=8'h00; mem['h2A7E]=8'h00; mem['h2A7F]=8'h00;
    mem['h2A80]=8'h00; mem['h2A81]=8'h00; mem['h2A82]=8'h00; mem['h2A83]=8'h00;
    mem['h2A84]=8'h00; mem['h2A85]=8'h00; mem['h2A86]=8'h00; mem['h2A87]=8'h00;
    mem['h2A88]=8'h00; mem['h2A89]=8'h00; mem['h2A8A]=8'h00; mem['h2A8B]=8'h00;
    mem['h2A8C]=8'h00; mem['h2A8D]=8'h00; mem['h2A8E]=8'h00; mem['h2A8F]=8'h00;
    mem['h2A90]=8'h00; mem['h2A91]=8'h00; mem['h2A92]=8'h00; mem['h2A93]=8'h00;
    mem['h2A94]=8'h00; mem['h2A95]=8'h00; mem['h2A96]=8'h00; mem['h2A97]=8'h00;
    mem['h2A98]=8'h00; mem['h2A99]=8'h00; mem['h2A9A]=8'h00; mem['h2A9B]=8'h00;
    mem['h2A9C]=8'h00; mem['h2A9D]=8'h00; mem['h2A9E]=8'h00; mem['h2A9F]=8'h00;
    mem['h2AA0]=8'h00; mem['h2AA1]=8'h00; mem['h2AA2]=8'h00; mem['h2AA3]=8'h00;
    mem['h2AA4]=8'h00; mem['h2AA5]=8'h00; mem['h2AA6]=8'h00; mem['h2AA7]=8'h00;
    mem['h2AA8]=8'h00; mem['h2AA9]=8'h00; mem['h2AAA]=8'h00; mem['h2AAB]=8'h00;
    mem['h2AAC]=8'h00; mem['h2AAD]=8'h00; mem['h2AAE]=8'h00; mem['h2AAF]=8'h00;
    mem['h2AB0]=8'h00; mem['h2AB1]=8'h00; mem['h2AB2]=8'h00; mem['h2AB3]=8'h00;
    mem['h2AB4]=8'h00; mem['h2AB5]=8'h00; mem['h2AB6]=8'h00; mem['h2AB7]=8'h00;
    mem['h2AB8]=8'h00; mem['h2AB9]=8'h00; mem['h2ABA]=8'h00; mem['h2ABB]=8'h00;
    mem['h2ABC]=8'h00; mem['h2ABD]=8'h00; mem['h2ABE]=8'h00; mem['h2ABF]=8'h00;
    mem['h2AC0]=8'h00; mem['h2AC1]=8'h00; mem['h2AC2]=8'h00; mem['h2AC3]=8'h00;
    mem['h2AC4]=8'h00; mem['h2AC5]=8'h00; mem['h2AC6]=8'h00; mem['h2AC7]=8'h00;
    mem['h2AC8]=8'h00; mem['h2AC9]=8'h00; mem['h2ACA]=8'h00; mem['h2ACB]=8'h00;
    mem['h2ACC]=8'h00; mem['h2ACD]=8'h00; mem['h2ACE]=8'h00; mem['h2ACF]=8'h00;
    mem['h2AD0]=8'h00; mem['h2AD1]=8'h00; mem['h2AD2]=8'h00; mem['h2AD3]=8'h00;
    mem['h2AD4]=8'h00; mem['h2AD5]=8'h00; mem['h2AD6]=8'h00; mem['h2AD7]=8'h00;
    mem['h2AD8]=8'h00; mem['h2AD9]=8'h00; mem['h2ADA]=8'h00; mem['h2ADB]=8'h00;
    mem['h2ADC]=8'h00; mem['h2ADD]=8'h00; mem['h2ADE]=8'h00; mem['h2ADF]=8'h00;
    mem['h2AE0]=8'h00; mem['h2AE1]=8'h00; mem['h2AE2]=8'h00; mem['h2AE3]=8'h00;
    mem['h2AE4]=8'h00; mem['h2AE5]=8'h00; mem['h2AE6]=8'h00; mem['h2AE7]=8'h00;
    mem['h2AE8]=8'h00; mem['h2AE9]=8'h00; mem['h2AEA]=8'h00; mem['h2AEB]=8'h00;
    mem['h2AEC]=8'h00; mem['h2AED]=8'h00; mem['h2AEE]=8'h00; mem['h2AEF]=8'h00;
    mem['h2AF0]=8'h00; mem['h2AF1]=8'h00; mem['h2AF2]=8'h00; mem['h2AF3]=8'h00;
    mem['h2AF4]=8'h00; mem['h2AF5]=8'h00; mem['h2AF6]=8'h00; mem['h2AF7]=8'h00;
    mem['h2AF8]=8'h00; mem['h2AF9]=8'h00; mem['h2AFA]=8'h00; mem['h2AFB]=8'h00;
    mem['h2AFC]=8'h00; mem['h2AFD]=8'h00; mem['h2AFE]=8'h00; mem['h2AFF]=8'h00;
    mem['h2B00]=8'h00; mem['h2B01]=8'h00; mem['h2B02]=8'h00; mem['h2B03]=8'h00;
    mem['h2B04]=8'h00; mem['h2B05]=8'h00; mem['h2B06]=8'h00; mem['h2B07]=8'h00;
    mem['h2B08]=8'h00; mem['h2B09]=8'h00; mem['h2B0A]=8'h00; mem['h2B0B]=8'h00;
    mem['h2B0C]=8'h00; mem['h2B0D]=8'h00; mem['h2B0E]=8'h00; mem['h2B0F]=8'h00;
    mem['h2B10]=8'h00; mem['h2B11]=8'h00; mem['h2B12]=8'h00; mem['h2B13]=8'h00;
    mem['h2B14]=8'h00; mem['h2B15]=8'h00; mem['h2B16]=8'h00; mem['h2B17]=8'h00;
    mem['h2B18]=8'h00; mem['h2B19]=8'h00; mem['h2B1A]=8'h00; mem['h2B1B]=8'h00;
    mem['h2B1C]=8'h00; mem['h2B1D]=8'h00; mem['h2B1E]=8'h00; mem['h2B1F]=8'h00;
    mem['h2B20]=8'h00; mem['h2B21]=8'h00; mem['h2B22]=8'h00; mem['h2B23]=8'h00;
    mem['h2B24]=8'h00; mem['h2B25]=8'h00; mem['h2B26]=8'h00; mem['h2B27]=8'h00;
    mem['h2B28]=8'h00; mem['h2B29]=8'h00; mem['h2B2A]=8'h00; mem['h2B2B]=8'h00;
    mem['h2B2C]=8'h00; mem['h2B2D]=8'h00; mem['h2B2E]=8'h00; mem['h2B2F]=8'h00;
    mem['h2B30]=8'h00; mem['h2B31]=8'h00; mem['h2B32]=8'h00; mem['h2B33]=8'h00;
    mem['h2B34]=8'h00; mem['h2B35]=8'h00; mem['h2B36]=8'h00; mem['h2B37]=8'h00;
    mem['h2B38]=8'h00; mem['h2B39]=8'h00; mem['h2B3A]=8'h00; mem['h2B3B]=8'h00;
    mem['h2B3C]=8'h00; mem['h2B3D]=8'h00; mem['h2B3E]=8'h00; mem['h2B3F]=8'h00;
    mem['h2B40]=8'h00; mem['h2B41]=8'h00; mem['h2B42]=8'h00; mem['h2B43]=8'h00;
    mem['h2B44]=8'h00; mem['h2B45]=8'h00; mem['h2B46]=8'h00; mem['h2B47]=8'h00;
    mem['h2B48]=8'h00; mem['h2B49]=8'h00; mem['h2B4A]=8'h00; mem['h2B4B]=8'h00;
    mem['h2B4C]=8'h00; mem['h2B4D]=8'h00; mem['h2B4E]=8'h00; mem['h2B4F]=8'h00;
    mem['h2B50]=8'h00; mem['h2B51]=8'h00; mem['h2B52]=8'h00; mem['h2B53]=8'h00;
    mem['h2B54]=8'h00; mem['h2B55]=8'h00; mem['h2B56]=8'h00; mem['h2B57]=8'h00;
    mem['h2B58]=8'h00; mem['h2B59]=8'h00; mem['h2B5A]=8'h00; mem['h2B5B]=8'h00;
    mem['h2B5C]=8'h00; mem['h2B5D]=8'h00; mem['h2B5E]=8'h00; mem['h2B5F]=8'h00;
    mem['h2B60]=8'h00; mem['h2B61]=8'h00; mem['h2B62]=8'h00; mem['h2B63]=8'h00;
    mem['h2B64]=8'h00; mem['h2B65]=8'h00; mem['h2B66]=8'h00; mem['h2B67]=8'h00;
    mem['h2B68]=8'h00; mem['h2B69]=8'h00; mem['h2B6A]=8'h00; mem['h2B6B]=8'h00;
    mem['h2B6C]=8'h00; mem['h2B6D]=8'h00; mem['h2B6E]=8'h00; mem['h2B6F]=8'h00;
    mem['h2B70]=8'h00; mem['h2B71]=8'h00; mem['h2B72]=8'h00; mem['h2B73]=8'h00;
    mem['h2B74]=8'h00; mem['h2B75]=8'h00; mem['h2B76]=8'h00; mem['h2B77]=8'h00;
    mem['h2B78]=8'h00; mem['h2B79]=8'h00; mem['h2B7A]=8'h00; mem['h2B7B]=8'h00;
    mem['h2B7C]=8'h00; mem['h2B7D]=8'h00; mem['h2B7E]=8'h00; mem['h2B7F]=8'h00;
    mem['h2B80]=8'h00; mem['h2B81]=8'h00; mem['h2B82]=8'h00; mem['h2B83]=8'h00;
    mem['h2B84]=8'h00; mem['h2B85]=8'h00; mem['h2B86]=8'h00; mem['h2B87]=8'h00;
    mem['h2B88]=8'h00; mem['h2B89]=8'h00; mem['h2B8A]=8'h00; mem['h2B8B]=8'h00;
    mem['h2B8C]=8'h00; mem['h2B8D]=8'h00; mem['h2B8E]=8'h00; mem['h2B8F]=8'h00;
    mem['h2B90]=8'h00; mem['h2B91]=8'h00; mem['h2B92]=8'h00; mem['h2B93]=8'h00;
    mem['h2B94]=8'h00; mem['h2B95]=8'h00; mem['h2B96]=8'h00; mem['h2B97]=8'h00;
    mem['h2B98]=8'h00; mem['h2B99]=8'h00; mem['h2B9A]=8'h00; mem['h2B9B]=8'h00;
    mem['h2B9C]=8'h00; mem['h2B9D]=8'h00; mem['h2B9E]=8'h00; mem['h2B9F]=8'h00;
    mem['h2BA0]=8'h00; mem['h2BA1]=8'h00; mem['h2BA2]=8'h00; mem['h2BA3]=8'h00;
    mem['h2BA4]=8'h00; mem['h2BA5]=8'h00; mem['h2BA6]=8'h00; mem['h2BA7]=8'h00;
    mem['h2BA8]=8'h00; mem['h2BA9]=8'h00; mem['h2BAA]=8'h00; mem['h2BAB]=8'h00;
    mem['h2BAC]=8'h00; mem['h2BAD]=8'h00; mem['h2BAE]=8'h00; mem['h2BAF]=8'h00;
    mem['h2BB0]=8'h00; mem['h2BB1]=8'h00; mem['h2BB2]=8'h00; mem['h2BB3]=8'h00;
    mem['h2BB4]=8'h00; mem['h2BB5]=8'h00; mem['h2BB6]=8'h00; mem['h2BB7]=8'h00;
    mem['h2BB8]=8'h00; mem['h2BB9]=8'h00; mem['h2BBA]=8'h00; mem['h2BBB]=8'h00;
    mem['h2BBC]=8'h00; mem['h2BBD]=8'h00; mem['h2BBE]=8'h00; mem['h2BBF]=8'h00;
    mem['h2BC0]=8'h00; mem['h2BC1]=8'h00; mem['h2BC2]=8'h00; mem['h2BC3]=8'h00;
    mem['h2BC4]=8'h00; mem['h2BC5]=8'h00; mem['h2BC6]=8'h00; mem['h2BC7]=8'h00;
    mem['h2BC8]=8'h00; mem['h2BC9]=8'h00; mem['h2BCA]=8'h00; mem['h2BCB]=8'h00;
    mem['h2BCC]=8'h00; mem['h2BCD]=8'h00; mem['h2BCE]=8'h00; mem['h2BCF]=8'h00;
    mem['h2BD0]=8'h00; mem['h2BD1]=8'h00; mem['h2BD2]=8'h00; mem['h2BD3]=8'h00;
    mem['h2BD4]=8'h00; mem['h2BD5]=8'h00; mem['h2BD6]=8'h00; mem['h2BD7]=8'h00;
    mem['h2BD8]=8'h00; mem['h2BD9]=8'h00; mem['h2BDA]=8'h00; mem['h2BDB]=8'h00;
    mem['h2BDC]=8'h00; mem['h2BDD]=8'h00; mem['h2BDE]=8'h00; mem['h2BDF]=8'h00;
    mem['h2BE0]=8'h00; mem['h2BE1]=8'h00; mem['h2BE2]=8'h00; mem['h2BE3]=8'h00;
    mem['h2BE4]=8'h00; mem['h2BE5]=8'h00; mem['h2BE6]=8'h00; mem['h2BE7]=8'h00;
    mem['h2BE8]=8'h00; mem['h2BE9]=8'h00; mem['h2BEA]=8'h00; mem['h2BEB]=8'h00;
    mem['h2BEC]=8'h00; mem['h2BED]=8'h00; mem['h2BEE]=8'h00; mem['h2BEF]=8'h00;
    mem['h2BF0]=8'h00; mem['h2BF1]=8'h00; mem['h2BF2]=8'h00; mem['h2BF3]=8'h00;
    mem['h2BF4]=8'h00; mem['h2BF5]=8'h00; mem['h2BF6]=8'h00; mem['h2BF7]=8'h00;
    mem['h2BF8]=8'h00; mem['h2BF9]=8'h00; mem['h2BFA]=8'h00; mem['h2BFB]=8'h00;
    mem['h2BFC]=8'h00; mem['h2BFD]=8'h00; mem['h2BFE]=8'h00; mem['h2BFF]=8'h00;
    mem['h2C00]=8'h00; mem['h2C01]=8'h00; mem['h2C02]=8'h00; mem['h2C03]=8'h00;
    mem['h2C04]=8'h00; mem['h2C05]=8'h00; mem['h2C06]=8'h00; mem['h2C07]=8'h00;
    mem['h2C08]=8'h00; mem['h2C09]=8'h00; mem['h2C0A]=8'h00; mem['h2C0B]=8'h00;
    mem['h2C0C]=8'h00; mem['h2C0D]=8'h00; mem['h2C0E]=8'h00; mem['h2C0F]=8'h00;
    mem['h2C10]=8'h00; mem['h2C11]=8'h00; mem['h2C12]=8'h00; mem['h2C13]=8'h00;
    mem['h2C14]=8'h00; mem['h2C15]=8'h00; mem['h2C16]=8'h00; mem['h2C17]=8'h00;
    mem['h2C18]=8'h00; mem['h2C19]=8'h00; mem['h2C1A]=8'h00; mem['h2C1B]=8'h00;
    mem['h2C1C]=8'h00; mem['h2C1D]=8'h00; mem['h2C1E]=8'h00; mem['h2C1F]=8'h00;
    mem['h2C20]=8'h00; mem['h2C21]=8'h00; mem['h2C22]=8'h00; mem['h2C23]=8'h00;
    mem['h2C24]=8'h00; mem['h2C25]=8'h00; mem['h2C26]=8'h00; mem['h2C27]=8'h00;
    mem['h2C28]=8'h00; mem['h2C29]=8'h00; mem['h2C2A]=8'h00; mem['h2C2B]=8'h00;
    mem['h2C2C]=8'h00; mem['h2C2D]=8'h00; mem['h2C2E]=8'h00; mem['h2C2F]=8'h00;
    mem['h2C30]=8'h00; mem['h2C31]=8'h00; mem['h2C32]=8'h00; mem['h2C33]=8'h00;
    mem['h2C34]=8'h00; mem['h2C35]=8'h00; mem['h2C36]=8'h00; mem['h2C37]=8'h00;
    mem['h2C38]=8'h00; mem['h2C39]=8'h00; mem['h2C3A]=8'h00; mem['h2C3B]=8'h00;
    mem['h2C3C]=8'h00; mem['h2C3D]=8'h00; mem['h2C3E]=8'h00; mem['h2C3F]=8'h00;
    mem['h2C40]=8'h00; mem['h2C41]=8'h00; mem['h2C42]=8'h00; mem['h2C43]=8'h00;
    mem['h2C44]=8'h00; mem['h2C45]=8'h00; mem['h2C46]=8'h00; mem['h2C47]=8'h00;
    mem['h2C48]=8'h00; mem['h2C49]=8'h00; mem['h2C4A]=8'h00; mem['h2C4B]=8'h00;
    mem['h2C4C]=8'h00; mem['h2C4D]=8'h00; mem['h2C4E]=8'h00; mem['h2C4F]=8'h00;
    mem['h2C50]=8'h00; mem['h2C51]=8'h00; mem['h2C52]=8'h00; mem['h2C53]=8'h00;
    mem['h2C54]=8'h00; mem['h2C55]=8'h00; mem['h2C56]=8'h00; mem['h2C57]=8'h00;
    mem['h2C58]=8'h00; mem['h2C59]=8'h00; mem['h2C5A]=8'h00; mem['h2C5B]=8'h00;
    mem['h2C5C]=8'h00; mem['h2C5D]=8'h00; mem['h2C5E]=8'h00; mem['h2C5F]=8'h00;
    mem['h2C60]=8'h00; mem['h2C61]=8'h00; mem['h2C62]=8'h00; mem['h2C63]=8'h00;
    mem['h2C64]=8'h00; mem['h2C65]=8'h00; mem['h2C66]=8'h00; mem['h2C67]=8'h00;
    mem['h2C68]=8'h00; mem['h2C69]=8'h00; mem['h2C6A]=8'h00; mem['h2C6B]=8'h00;
    mem['h2C6C]=8'h00; mem['h2C6D]=8'h00; mem['h2C6E]=8'h00; mem['h2C6F]=8'h00;
    mem['h2C70]=8'h00; mem['h2C71]=8'h00; mem['h2C72]=8'h00; mem['h2C73]=8'h00;
    mem['h2C74]=8'h00; mem['h2C75]=8'h00; mem['h2C76]=8'h00; mem['h2C77]=8'h00;
    mem['h2C78]=8'h00; mem['h2C79]=8'h00; mem['h2C7A]=8'h00; mem['h2C7B]=8'h00;
    mem['h2C7C]=8'h00; mem['h2C7D]=8'h00; mem['h2C7E]=8'h00; mem['h2C7F]=8'h00;
    mem['h2C80]=8'h00; mem['h2C81]=8'h00; mem['h2C82]=8'h00; mem['h2C83]=8'h00;
    mem['h2C84]=8'h00; mem['h2C85]=8'h00; mem['h2C86]=8'h00; mem['h2C87]=8'h00;
    mem['h2C88]=8'h00; mem['h2C89]=8'h00; mem['h2C8A]=8'h00; mem['h2C8B]=8'h00;
    mem['h2C8C]=8'h00; mem['h2C8D]=8'h00; mem['h2C8E]=8'h00; mem['h2C8F]=8'h00;
    mem['h2C90]=8'h00; mem['h2C91]=8'h00; mem['h2C92]=8'h00; mem['h2C93]=8'h00;
    mem['h2C94]=8'h00; mem['h2C95]=8'h00; mem['h2C96]=8'h00; mem['h2C97]=8'h00;
    mem['h2C98]=8'h00; mem['h2C99]=8'h00; mem['h2C9A]=8'h00; mem['h2C9B]=8'h00;
    mem['h2C9C]=8'h00; mem['h2C9D]=8'h00; mem['h2C9E]=8'h00; mem['h2C9F]=8'h00;
    mem['h2CA0]=8'h00; mem['h2CA1]=8'h00; mem['h2CA2]=8'h00; mem['h2CA3]=8'h00;
    mem['h2CA4]=8'h00; mem['h2CA5]=8'h00; mem['h2CA6]=8'h00; mem['h2CA7]=8'h00;
    mem['h2CA8]=8'h00; mem['h2CA9]=8'h00; mem['h2CAA]=8'h00; mem['h2CAB]=8'h00;
    mem['h2CAC]=8'h00; mem['h2CAD]=8'h00; mem['h2CAE]=8'h00; mem['h2CAF]=8'h00;
    mem['h2CB0]=8'h00; mem['h2CB1]=8'h00; mem['h2CB2]=8'h00; mem['h2CB3]=8'h00;
    mem['h2CB4]=8'h00; mem['h2CB5]=8'h00; mem['h2CB6]=8'h00; mem['h2CB7]=8'h00;
    mem['h2CB8]=8'h00; mem['h2CB9]=8'h00; mem['h2CBA]=8'h00; mem['h2CBB]=8'h00;
    mem['h2CBC]=8'h00; mem['h2CBD]=8'h00; mem['h2CBE]=8'h00; mem['h2CBF]=8'h00;
    mem['h2CC0]=8'h00; mem['h2CC1]=8'h00; mem['h2CC2]=8'h00; mem['h2CC3]=8'h00;
    mem['h2CC4]=8'h00; mem['h2CC5]=8'h00; mem['h2CC6]=8'h00; mem['h2CC7]=8'h00;
    mem['h2CC8]=8'h00; mem['h2CC9]=8'h00; mem['h2CCA]=8'h00; mem['h2CCB]=8'h00;
    mem['h2CCC]=8'h00; mem['h2CCD]=8'h00; mem['h2CCE]=8'h00; mem['h2CCF]=8'h00;
    mem['h2CD0]=8'h00; mem['h2CD1]=8'h00; mem['h2CD2]=8'h00; mem['h2CD3]=8'h00;
    mem['h2CD4]=8'h00; mem['h2CD5]=8'h00; mem['h2CD6]=8'h00; mem['h2CD7]=8'h00;
    mem['h2CD8]=8'h00; mem['h2CD9]=8'h00; mem['h2CDA]=8'h00; mem['h2CDB]=8'h00;
    mem['h2CDC]=8'h00; mem['h2CDD]=8'h00; mem['h2CDE]=8'h00; mem['h2CDF]=8'h00;
    mem['h2CE0]=8'h00; mem['h2CE1]=8'h00; mem['h2CE2]=8'h00; mem['h2CE3]=8'h00;
    mem['h2CE4]=8'h00; mem['h2CE5]=8'h00; mem['h2CE6]=8'h00; mem['h2CE7]=8'h00;
    mem['h2CE8]=8'h00; mem['h2CE9]=8'h00; mem['h2CEA]=8'h00; mem['h2CEB]=8'h00;
    mem['h2CEC]=8'h00; mem['h2CED]=8'h00; mem['h2CEE]=8'h00; mem['h2CEF]=8'h00;
    mem['h2CF0]=8'h00; mem['h2CF1]=8'h00; mem['h2CF2]=8'h00; mem['h2CF3]=8'h00;
    mem['h2CF4]=8'h00; mem['h2CF5]=8'h00; mem['h2CF6]=8'h00; mem['h2CF7]=8'h00;
    mem['h2CF8]=8'h00; mem['h2CF9]=8'h00; mem['h2CFA]=8'h00; mem['h2CFB]=8'h00;
    mem['h2CFC]=8'h00; mem['h2CFD]=8'h00; mem['h2CFE]=8'h00; mem['h2CFF]=8'h00;
    mem['h2D00]=8'h00; mem['h2D01]=8'h00; mem['h2D02]=8'h00; mem['h2D03]=8'h00;
    mem['h2D04]=8'h00; mem['h2D05]=8'h00; mem['h2D06]=8'h00; mem['h2D07]=8'h00;
    mem['h2D08]=8'h00; mem['h2D09]=8'h00; mem['h2D0A]=8'h00; mem['h2D0B]=8'h00;
    mem['h2D0C]=8'h00; mem['h2D0D]=8'h00; mem['h2D0E]=8'h00; mem['h2D0F]=8'h00;
    mem['h2D10]=8'h00; mem['h2D11]=8'h00; mem['h2D12]=8'h00; mem['h2D13]=8'h00;
    mem['h2D14]=8'h00; mem['h2D15]=8'h00; mem['h2D16]=8'h00; mem['h2D17]=8'h00;
    mem['h2D18]=8'h00; mem['h2D19]=8'h00; mem['h2D1A]=8'h00; mem['h2D1B]=8'h00;
    mem['h2D1C]=8'h00; mem['h2D1D]=8'h00; mem['h2D1E]=8'h00; mem['h2D1F]=8'h00;
    mem['h2D20]=8'h00; mem['h2D21]=8'h00; mem['h2D22]=8'h00; mem['h2D23]=8'h00;
    mem['h2D24]=8'h00; mem['h2D25]=8'h00; mem['h2D26]=8'h00; mem['h2D27]=8'h00;
    mem['h2D28]=8'h00; mem['h2D29]=8'h00; mem['h2D2A]=8'h00; mem['h2D2B]=8'h00;
    mem['h2D2C]=8'h00; mem['h2D2D]=8'h00; mem['h2D2E]=8'h00; mem['h2D2F]=8'h00;
    mem['h2D30]=8'h00; mem['h2D31]=8'h00; mem['h2D32]=8'h00; mem['h2D33]=8'h00;
    mem['h2D34]=8'h00; mem['h2D35]=8'h00; mem['h2D36]=8'h00; mem['h2D37]=8'h00;
    mem['h2D38]=8'h00; mem['h2D39]=8'h00; mem['h2D3A]=8'h00; mem['h2D3B]=8'h00;
    mem['h2D3C]=8'h00; mem['h2D3D]=8'h00; mem['h2D3E]=8'h00; mem['h2D3F]=8'h00;
    mem['h2D40]=8'h00; mem['h2D41]=8'h00; mem['h2D42]=8'h00; mem['h2D43]=8'h00;
    mem['h2D44]=8'h00; mem['h2D45]=8'h00; mem['h2D46]=8'h00; mem['h2D47]=8'h00;
    mem['h2D48]=8'h00; mem['h2D49]=8'h00; mem['h2D4A]=8'h00; mem['h2D4B]=8'h00;
    mem['h2D4C]=8'h00; mem['h2D4D]=8'h00; mem['h2D4E]=8'h00; mem['h2D4F]=8'h00;
    mem['h2D50]=8'h00; mem['h2D51]=8'h00; mem['h2D52]=8'h00; mem['h2D53]=8'h00;
    mem['h2D54]=8'h00; mem['h2D55]=8'h00; mem['h2D56]=8'h00; mem['h2D57]=8'h00;
    mem['h2D58]=8'h00; mem['h2D59]=8'h00; mem['h2D5A]=8'h00; mem['h2D5B]=8'h00;
    mem['h2D5C]=8'h00; mem['h2D5D]=8'h00; mem['h2D5E]=8'h00; mem['h2D5F]=8'h00;
    mem['h2D60]=8'h00; mem['h2D61]=8'h00; mem['h2D62]=8'h00; mem['h2D63]=8'h00;
    mem['h2D64]=8'h00; mem['h2D65]=8'h00; mem['h2D66]=8'h00; mem['h2D67]=8'h00;
    mem['h2D68]=8'h00; mem['h2D69]=8'h00; mem['h2D6A]=8'h00; mem['h2D6B]=8'h00;
    mem['h2D6C]=8'h00; mem['h2D6D]=8'h00; mem['h2D6E]=8'h00; mem['h2D6F]=8'h00;
    mem['h2D70]=8'h00; mem['h2D71]=8'h00; mem['h2D72]=8'h00; mem['h2D73]=8'h00;
    mem['h2D74]=8'h00; mem['h2D75]=8'h00; mem['h2D76]=8'h00; mem['h2D77]=8'h00;
    mem['h2D78]=8'h00; mem['h2D79]=8'h00; mem['h2D7A]=8'h00; mem['h2D7B]=8'h00;
    mem['h2D7C]=8'h00; mem['h2D7D]=8'h00; mem['h2D7E]=8'h00; mem['h2D7F]=8'h00;
    mem['h2D80]=8'h00; mem['h2D81]=8'h00; mem['h2D82]=8'h00; mem['h2D83]=8'h00;
    mem['h2D84]=8'h00; mem['h2D85]=8'h00; mem['h2D86]=8'h00; mem['h2D87]=8'h00;
    mem['h2D88]=8'h00; mem['h2D89]=8'h00; mem['h2D8A]=8'h00; mem['h2D8B]=8'h00;
    mem['h2D8C]=8'h00; mem['h2D8D]=8'h00; mem['h2D8E]=8'h00; mem['h2D8F]=8'h00;
    mem['h2D90]=8'h00; mem['h2D91]=8'h00; mem['h2D92]=8'h00; mem['h2D93]=8'h00;
    mem['h2D94]=8'h00; mem['h2D95]=8'h00; mem['h2D96]=8'h00; mem['h2D97]=8'h00;
    mem['h2D98]=8'h00; mem['h2D99]=8'h00; mem['h2D9A]=8'h00; mem['h2D9B]=8'h00;
    mem['h2D9C]=8'h00; mem['h2D9D]=8'h00; mem['h2D9E]=8'h00; mem['h2D9F]=8'h00;
    mem['h2DA0]=8'h00; mem['h2DA1]=8'h00; mem['h2DA2]=8'h00; mem['h2DA3]=8'h00;
    mem['h2DA4]=8'h00; mem['h2DA5]=8'h00; mem['h2DA6]=8'h00; mem['h2DA7]=8'h00;
    mem['h2DA8]=8'h00; mem['h2DA9]=8'h00; mem['h2DAA]=8'h00; mem['h2DAB]=8'h00;
    mem['h2DAC]=8'h00; mem['h2DAD]=8'h00; mem['h2DAE]=8'h00; mem['h2DAF]=8'h00;
    mem['h2DB0]=8'h00; mem['h2DB1]=8'h00; mem['h2DB2]=8'h00; mem['h2DB3]=8'h00;
    mem['h2DB4]=8'h00; mem['h2DB5]=8'h00; mem['h2DB6]=8'h00; mem['h2DB7]=8'h00;
    mem['h2DB8]=8'h00; mem['h2DB9]=8'h00; mem['h2DBA]=8'h00; mem['h2DBB]=8'h00;
    mem['h2DBC]=8'h00; mem['h2DBD]=8'h00; mem['h2DBE]=8'h00; mem['h2DBF]=8'h00;
    mem['h2DC0]=8'h00; mem['h2DC1]=8'h00; mem['h2DC2]=8'h00; mem['h2DC3]=8'h00;
    mem['h2DC4]=8'h00; mem['h2DC5]=8'h00; mem['h2DC6]=8'h00; mem['h2DC7]=8'h00;
    mem['h2DC8]=8'h00; mem['h2DC9]=8'h00; mem['h2DCA]=8'h00; mem['h2DCB]=8'h00;
    mem['h2DCC]=8'h00; mem['h2DCD]=8'h00; mem['h2DCE]=8'h00; mem['h2DCF]=8'h00;
    mem['h2DD0]=8'h00; mem['h2DD1]=8'h00; mem['h2DD2]=8'h00; mem['h2DD3]=8'h00;
    mem['h2DD4]=8'h00; mem['h2DD5]=8'h00; mem['h2DD6]=8'h00; mem['h2DD7]=8'h00;
    mem['h2DD8]=8'h00; mem['h2DD9]=8'h00; mem['h2DDA]=8'h00; mem['h2DDB]=8'h00;
    mem['h2DDC]=8'h00; mem['h2DDD]=8'h00; mem['h2DDE]=8'h00; mem['h2DDF]=8'h00;
    mem['h2DE0]=8'h00; mem['h2DE1]=8'h00; mem['h2DE2]=8'h00; mem['h2DE3]=8'h00;
    mem['h2DE4]=8'h00; mem['h2DE5]=8'h00; mem['h2DE6]=8'h00; mem['h2DE7]=8'h00;
    mem['h2DE8]=8'h00; mem['h2DE9]=8'h00; mem['h2DEA]=8'h00; mem['h2DEB]=8'h00;
    mem['h2DEC]=8'h00; mem['h2DED]=8'h00; mem['h2DEE]=8'h00; mem['h2DEF]=8'h00;
    mem['h2DF0]=8'h00; mem['h2DF1]=8'h00; mem['h2DF2]=8'h00; mem['h2DF3]=8'h00;
    mem['h2DF4]=8'h00; mem['h2DF5]=8'h00; mem['h2DF6]=8'h00; mem['h2DF7]=8'h00;
    mem['h2DF8]=8'h00; mem['h2DF9]=8'h00; mem['h2DFA]=8'h00; mem['h2DFB]=8'h00;
    mem['h2DFC]=8'h00; mem['h2DFD]=8'h00; mem['h2DFE]=8'h00; mem['h2DFF]=8'h00;
    mem['h2E00]=8'h00; mem['h2E01]=8'h00; mem['h2E02]=8'h00; mem['h2E03]=8'h00;
    mem['h2E04]=8'h00; mem['h2E05]=8'h00; mem['h2E06]=8'h00; mem['h2E07]=8'h00;
    mem['h2E08]=8'h00; mem['h2E09]=8'h00; mem['h2E0A]=8'h00; mem['h2E0B]=8'h00;
    mem['h2E0C]=8'h00; mem['h2E0D]=8'h00; mem['h2E0E]=8'h00; mem['h2E0F]=8'h00;
    mem['h2E10]=8'h00; mem['h2E11]=8'h00; mem['h2E12]=8'h00; mem['h2E13]=8'h00;
    mem['h2E14]=8'h00; mem['h2E15]=8'h00; mem['h2E16]=8'h00; mem['h2E17]=8'h00;
    mem['h2E18]=8'h00; mem['h2E19]=8'h00; mem['h2E1A]=8'h00; mem['h2E1B]=8'h00;
    mem['h2E1C]=8'h00; mem['h2E1D]=8'h00; mem['h2E1E]=8'h00; mem['h2E1F]=8'h00;
    mem['h2E20]=8'h00; mem['h2E21]=8'h00; mem['h2E22]=8'h00; mem['h2E23]=8'h00;
    mem['h2E24]=8'h00; mem['h2E25]=8'h00; mem['h2E26]=8'h00; mem['h2E27]=8'h00;
    mem['h2E28]=8'h00; mem['h2E29]=8'h00; mem['h2E2A]=8'h00; mem['h2E2B]=8'h00;
    mem['h2E2C]=8'h00; mem['h2E2D]=8'h00; mem['h2E2E]=8'h00; mem['h2E2F]=8'h00;
    mem['h2E30]=8'h00; mem['h2E31]=8'h00; mem['h2E32]=8'h00; mem['h2E33]=8'h00;
    mem['h2E34]=8'h00; mem['h2E35]=8'h00; mem['h2E36]=8'h00; mem['h2E37]=8'h00;
    mem['h2E38]=8'h00; mem['h2E39]=8'h00; mem['h2E3A]=8'h00; mem['h2E3B]=8'h00;
    mem['h2E3C]=8'h00; mem['h2E3D]=8'h00; mem['h2E3E]=8'h00; mem['h2E3F]=8'h00;
    mem['h2E40]=8'h00; mem['h2E41]=8'h00; mem['h2E42]=8'h00; mem['h2E43]=8'h00;
    mem['h2E44]=8'h00; mem['h2E45]=8'h00; mem['h2E46]=8'h00; mem['h2E47]=8'h00;
    mem['h2E48]=8'h00; mem['h2E49]=8'h00; mem['h2E4A]=8'h00; mem['h2E4B]=8'h00;
    mem['h2E4C]=8'h00; mem['h2E4D]=8'h00; mem['h2E4E]=8'h00; mem['h2E4F]=8'h00;
    mem['h2E50]=8'h00; mem['h2E51]=8'h00; mem['h2E52]=8'h00; mem['h2E53]=8'h00;
    mem['h2E54]=8'h00; mem['h2E55]=8'h00; mem['h2E56]=8'h00; mem['h2E57]=8'h00;
    mem['h2E58]=8'h00; mem['h2E59]=8'h00; mem['h2E5A]=8'h00; mem['h2E5B]=8'h00;
    mem['h2E5C]=8'h00; mem['h2E5D]=8'h00; mem['h2E5E]=8'h00; mem['h2E5F]=8'h00;
    mem['h2E60]=8'h00; mem['h2E61]=8'h00; mem['h2E62]=8'h00; mem['h2E63]=8'h00;
    mem['h2E64]=8'h00; mem['h2E65]=8'h00; mem['h2E66]=8'h00; mem['h2E67]=8'h00;
    mem['h2E68]=8'h00; mem['h2E69]=8'h00; mem['h2E6A]=8'h00; mem['h2E6B]=8'h00;
    mem['h2E6C]=8'h00; mem['h2E6D]=8'h00; mem['h2E6E]=8'h00; mem['h2E6F]=8'h00;
    mem['h2E70]=8'h00; mem['h2E71]=8'h00; mem['h2E72]=8'h00; mem['h2E73]=8'h00;
    mem['h2E74]=8'h00; mem['h2E75]=8'h00; mem['h2E76]=8'h00; mem['h2E77]=8'h00;
    mem['h2E78]=8'h00; mem['h2E79]=8'h00; mem['h2E7A]=8'h00; mem['h2E7B]=8'h00;
    mem['h2E7C]=8'h00; mem['h2E7D]=8'h00; mem['h2E7E]=8'h00; mem['h2E7F]=8'h00;
    mem['h2E80]=8'h00; mem['h2E81]=8'h00; mem['h2E82]=8'h00; mem['h2E83]=8'h00;
    mem['h2E84]=8'h00; mem['h2E85]=8'h00; mem['h2E86]=8'h00; mem['h2E87]=8'h00;
    mem['h2E88]=8'h00; mem['h2E89]=8'h00; mem['h2E8A]=8'h00; mem['h2E8B]=8'h00;
    mem['h2E8C]=8'h00; mem['h2E8D]=8'h00; mem['h2E8E]=8'h00; mem['h2E8F]=8'h00;
    mem['h2E90]=8'h00; mem['h2E91]=8'h00; mem['h2E92]=8'h00; mem['h2E93]=8'h00;
    mem['h2E94]=8'h00; mem['h2E95]=8'h00; mem['h2E96]=8'h00; mem['h2E97]=8'h00;
    mem['h2E98]=8'h00; mem['h2E99]=8'h00; mem['h2E9A]=8'h00; mem['h2E9B]=8'h00;
    mem['h2E9C]=8'h00; mem['h2E9D]=8'h00; mem['h2E9E]=8'h00; mem['h2E9F]=8'h00;
    mem['h2EA0]=8'h00; mem['h2EA1]=8'h00; mem['h2EA2]=8'h00; mem['h2EA3]=8'h00;
    mem['h2EA4]=8'h00; mem['h2EA5]=8'h00; mem['h2EA6]=8'h00; mem['h2EA7]=8'h00;
    mem['h2EA8]=8'h00; mem['h2EA9]=8'h00; mem['h2EAA]=8'h00; mem['h2EAB]=8'h00;
    mem['h2EAC]=8'h00; mem['h2EAD]=8'h00; mem['h2EAE]=8'h00; mem['h2EAF]=8'h00;
    mem['h2EB0]=8'h00; mem['h2EB1]=8'h00; mem['h2EB2]=8'h00; mem['h2EB3]=8'h00;
    mem['h2EB4]=8'h00; mem['h2EB5]=8'h00; mem['h2EB6]=8'h00; mem['h2EB7]=8'h00;
    mem['h2EB8]=8'h00; mem['h2EB9]=8'h00; mem['h2EBA]=8'h00; mem['h2EBB]=8'h00;
    mem['h2EBC]=8'h00; mem['h2EBD]=8'h00; mem['h2EBE]=8'h00; mem['h2EBF]=8'h00;
    mem['h2EC0]=8'h00; mem['h2EC1]=8'h00; mem['h2EC2]=8'h00; mem['h2EC3]=8'h00;
    mem['h2EC4]=8'h00; mem['h2EC5]=8'h00; mem['h2EC6]=8'h00; mem['h2EC7]=8'h00;
    mem['h2EC8]=8'h00; mem['h2EC9]=8'h00; mem['h2ECA]=8'h00; mem['h2ECB]=8'h00;
    mem['h2ECC]=8'h00; mem['h2ECD]=8'h00; mem['h2ECE]=8'h00; mem['h2ECF]=8'h00;
    mem['h2ED0]=8'h00; mem['h2ED1]=8'h00; mem['h2ED2]=8'h00; mem['h2ED3]=8'h00;
    mem['h2ED4]=8'h00; mem['h2ED5]=8'h00; mem['h2ED6]=8'h00; mem['h2ED7]=8'h00;
    mem['h2ED8]=8'h00; mem['h2ED9]=8'h00; mem['h2EDA]=8'h00; mem['h2EDB]=8'h00;
    mem['h2EDC]=8'h00; mem['h2EDD]=8'h00; mem['h2EDE]=8'h00; mem['h2EDF]=8'h00;
    mem['h2EE0]=8'h00; mem['h2EE1]=8'h00; mem['h2EE2]=8'h00; mem['h2EE3]=8'h00;
    mem['h2EE4]=8'h00; mem['h2EE5]=8'h00; mem['h2EE6]=8'h00; mem['h2EE7]=8'h00;
    mem['h2EE8]=8'h00; mem['h2EE9]=8'h00; mem['h2EEA]=8'h00; mem['h2EEB]=8'h00;
    mem['h2EEC]=8'h00; mem['h2EED]=8'h00; mem['h2EEE]=8'h00; mem['h2EEF]=8'h00;
    mem['h2EF0]=8'h00; mem['h2EF1]=8'h00; mem['h2EF2]=8'h00; mem['h2EF3]=8'h00;
    mem['h2EF4]=8'h00; mem['h2EF5]=8'h00; mem['h2EF6]=8'h00; mem['h2EF7]=8'h00;
    mem['h2EF8]=8'h00; mem['h2EF9]=8'h00; mem['h2EFA]=8'h00; mem['h2EFB]=8'h00;
    mem['h2EFC]=8'h00; mem['h2EFD]=8'h00; mem['h2EFE]=8'h00; mem['h2EFF]=8'h00;
    mem['h2F00]=8'h00; mem['h2F01]=8'h00; mem['h2F02]=8'h00; mem['h2F03]=8'h00;
    mem['h2F04]=8'h00; mem['h2F05]=8'h00; mem['h2F06]=8'h00; mem['h2F07]=8'h00;
    mem['h2F08]=8'h00; mem['h2F09]=8'h00; mem['h2F0A]=8'h00; mem['h2F0B]=8'h00;
    mem['h2F0C]=8'h00; mem['h2F0D]=8'h00; mem['h2F0E]=8'h00; mem['h2F0F]=8'h00;
    mem['h2F10]=8'h00; mem['h2F11]=8'h00; mem['h2F12]=8'h00; mem['h2F13]=8'h00;
    mem['h2F14]=8'h00; mem['h2F15]=8'h00; mem['h2F16]=8'h00; mem['h2F17]=8'h00;
    mem['h2F18]=8'h00; mem['h2F19]=8'h00; mem['h2F1A]=8'h00; mem['h2F1B]=8'h00;
    mem['h2F1C]=8'h00; mem['h2F1D]=8'h00; mem['h2F1E]=8'h00; mem['h2F1F]=8'h00;
    mem['h2F20]=8'h00; mem['h2F21]=8'h00; mem['h2F22]=8'h00; mem['h2F23]=8'h00;
    mem['h2F24]=8'h00; mem['h2F25]=8'h00; mem['h2F26]=8'h00; mem['h2F27]=8'h00;
    mem['h2F28]=8'h00; mem['h2F29]=8'h00; mem['h2F2A]=8'h00; mem['h2F2B]=8'h00;
    mem['h2F2C]=8'h00; mem['h2F2D]=8'h00; mem['h2F2E]=8'h00; mem['h2F2F]=8'h00;
    mem['h2F30]=8'h00; mem['h2F31]=8'h00; mem['h2F32]=8'h00; mem['h2F33]=8'h00;
    mem['h2F34]=8'h00; mem['h2F35]=8'h00; mem['h2F36]=8'h00; mem['h2F37]=8'h00;
    mem['h2F38]=8'h00; mem['h2F39]=8'h00; mem['h2F3A]=8'h00; mem['h2F3B]=8'h00;
    mem['h2F3C]=8'h00; mem['h2F3D]=8'h00; mem['h2F3E]=8'h00; mem['h2F3F]=8'h00;
    mem['h2F40]=8'h00; mem['h2F41]=8'h00; mem['h2F42]=8'h00; mem['h2F43]=8'h00;
    mem['h2F44]=8'h00; mem['h2F45]=8'h00; mem['h2F46]=8'h00; mem['h2F47]=8'h00;
    mem['h2F48]=8'h00; mem['h2F49]=8'h00; mem['h2F4A]=8'h00; mem['h2F4B]=8'h00;
    mem['h2F4C]=8'h00; mem['h2F4D]=8'h00; mem['h2F4E]=8'h00; mem['h2F4F]=8'h00;
    mem['h2F50]=8'h00; mem['h2F51]=8'h00; mem['h2F52]=8'h00; mem['h2F53]=8'h00;
    mem['h2F54]=8'h00; mem['h2F55]=8'h00; mem['h2F56]=8'h00; mem['h2F57]=8'h00;
    mem['h2F58]=8'h00; mem['h2F59]=8'h00; mem['h2F5A]=8'h00; mem['h2F5B]=8'h00;
    mem['h2F5C]=8'h00; mem['h2F5D]=8'h00; mem['h2F5E]=8'h00; mem['h2F5F]=8'h00;
    mem['h2F60]=8'h00; mem['h2F61]=8'h00; mem['h2F62]=8'h00; mem['h2F63]=8'h00;
    mem['h2F64]=8'h00; mem['h2F65]=8'h00; mem['h2F66]=8'h00; mem['h2F67]=8'h00;
    mem['h2F68]=8'h00; mem['h2F69]=8'h00; mem['h2F6A]=8'h00; mem['h2F6B]=8'h00;
    mem['h2F6C]=8'h00; mem['h2F6D]=8'h00; mem['h2F6E]=8'h00; mem['h2F6F]=8'h00;
    mem['h2F70]=8'h00; mem['h2F71]=8'h00; mem['h2F72]=8'h00; mem['h2F73]=8'h00;
    mem['h2F74]=8'h00; mem['h2F75]=8'h00; mem['h2F76]=8'h00; mem['h2F77]=8'h00;
    mem['h2F78]=8'h00; mem['h2F79]=8'h00; mem['h2F7A]=8'h00; mem['h2F7B]=8'h00;
    mem['h2F7C]=8'h00; mem['h2F7D]=8'h00; mem['h2F7E]=8'h00; mem['h2F7F]=8'h00;
    mem['h2F80]=8'h00; mem['h2F81]=8'h00; mem['h2F82]=8'h00; mem['h2F83]=8'h00;
    mem['h2F84]=8'h00; mem['h2F85]=8'h00; mem['h2F86]=8'h00; mem['h2F87]=8'h00;
    mem['h2F88]=8'h00; mem['h2F89]=8'h00; mem['h2F8A]=8'h00; mem['h2F8B]=8'h00;
    mem['h2F8C]=8'h00; mem['h2F8D]=8'h00; mem['h2F8E]=8'h00; mem['h2F8F]=8'h00;
    mem['h2F90]=8'h00; mem['h2F91]=8'h00; mem['h2F92]=8'h00; mem['h2F93]=8'h00;
    mem['h2F94]=8'h00; mem['h2F95]=8'h00; mem['h2F96]=8'h00; mem['h2F97]=8'h00;
    mem['h2F98]=8'h00; mem['h2F99]=8'h00; mem['h2F9A]=8'h00; mem['h2F9B]=8'h00;
    mem['h2F9C]=8'h00; mem['h2F9D]=8'h00; mem['h2F9E]=8'h00; mem['h2F9F]=8'h00;
    mem['h2FA0]=8'h00; mem['h2FA1]=8'h00; mem['h2FA2]=8'h00; mem['h2FA3]=8'h00;
    mem['h2FA4]=8'h00; mem['h2FA5]=8'h00; mem['h2FA6]=8'h00; mem['h2FA7]=8'h00;
    mem['h2FA8]=8'h00; mem['h2FA9]=8'h00; mem['h2FAA]=8'h00; mem['h2FAB]=8'h00;
    mem['h2FAC]=8'h00; mem['h2FAD]=8'h00; mem['h2FAE]=8'h00; mem['h2FAF]=8'h00;
    mem['h2FB0]=8'h00; mem['h2FB1]=8'h00; mem['h2FB2]=8'h00; mem['h2FB3]=8'h00;
    mem['h2FB4]=8'h00; mem['h2FB5]=8'h00; mem['h2FB6]=8'h00; mem['h2FB7]=8'h00;
    mem['h2FB8]=8'h00; mem['h2FB9]=8'h00; mem['h2FBA]=8'h00; mem['h2FBB]=8'h00;
    mem['h2FBC]=8'h00; mem['h2FBD]=8'h00; mem['h2FBE]=8'h00; mem['h2FBF]=8'h00;
    mem['h2FC0]=8'h00; mem['h2FC1]=8'h00; mem['h2FC2]=8'h00; mem['h2FC3]=8'h00;
    mem['h2FC4]=8'h00; mem['h2FC5]=8'h00; mem['h2FC6]=8'h00; mem['h2FC7]=8'h00;
    mem['h2FC8]=8'h00; mem['h2FC9]=8'h00; mem['h2FCA]=8'h00; mem['h2FCB]=8'h00;
    mem['h2FCC]=8'h00; mem['h2FCD]=8'h00; mem['h2FCE]=8'h00; mem['h2FCF]=8'h00;
    mem['h2FD0]=8'h00; mem['h2FD1]=8'h00; mem['h2FD2]=8'h00; mem['h2FD3]=8'h00;
    mem['h2FD4]=8'h00; mem['h2FD5]=8'h00; mem['h2FD6]=8'h00; mem['h2FD7]=8'h00;
    mem['h2FD8]=8'h00; mem['h2FD9]=8'h00; mem['h2FDA]=8'h00; mem['h2FDB]=8'h00;
    mem['h2FDC]=8'h00; mem['h2FDD]=8'h00; mem['h2FDE]=8'h00; mem['h2FDF]=8'h00;
    mem['h2FE0]=8'h00; mem['h2FE1]=8'h00; mem['h2FE2]=8'h00; mem['h2FE3]=8'h00;
    mem['h2FE4]=8'h00; mem['h2FE5]=8'h00; mem['h2FE6]=8'h00; mem['h2FE7]=8'h00;
    mem['h2FE8]=8'h00; mem['h2FE9]=8'h00; mem['h2FEA]=8'h00; mem['h2FEB]=8'h00;
    mem['h2FEC]=8'h00; mem['h2FED]=8'h00; mem['h2FEE]=8'h00; mem['h2FEF]=8'h00;
    mem['h2FF0]=8'h00; mem['h2FF1]=8'h00; mem['h2FF2]=8'h00; mem['h2FF3]=8'h00;
    mem['h2FF4]=8'h00; mem['h2FF5]=8'h00; mem['h2FF6]=8'h00; mem['h2FF7]=8'h00;
    mem['h2FF8]=8'h00; mem['h2FF9]=8'h00; mem['h2FFA]=8'h00; mem['h2FFB]=8'h00;
    mem['h2FFC]=8'h00; mem['h2FFD]=8'h00; mem['h2FFE]=8'h00; mem['h2FFF]=8'h00;
    mem['h3000]=8'h00; mem['h3001]=8'h00; mem['h3002]=8'h00; mem['h3003]=8'h00;
    mem['h3004]=8'h00; mem['h3005]=8'h00; mem['h3006]=8'h00; mem['h3007]=8'h00;
    mem['h3008]=8'h00; mem['h3009]=8'h00; mem['h300A]=8'h00; mem['h300B]=8'h00;
    mem['h300C]=8'h00; mem['h300D]=8'h00; mem['h300E]=8'h00; mem['h300F]=8'h00;
    mem['h3010]=8'h00; mem['h3011]=8'h00; mem['h3012]=8'h00; mem['h3013]=8'h00;
    mem['h3014]=8'h00; mem['h3015]=8'h00; mem['h3016]=8'h00; mem['h3017]=8'h00;
    mem['h3018]=8'h00; mem['h3019]=8'h00; mem['h301A]=8'h00; mem['h301B]=8'h00;
    mem['h301C]=8'h00; mem['h301D]=8'h00; mem['h301E]=8'h00; mem['h301F]=8'h00;
    mem['h3020]=8'h00; mem['h3021]=8'h00; mem['h3022]=8'h00; mem['h3023]=8'h00;
    mem['h3024]=8'h00; mem['h3025]=8'h00; mem['h3026]=8'h00; mem['h3027]=8'h00;
    mem['h3028]=8'h00; mem['h3029]=8'h00; mem['h302A]=8'h00; mem['h302B]=8'h00;
    mem['h302C]=8'h00; mem['h302D]=8'h00; mem['h302E]=8'h00; mem['h302F]=8'h00;
    mem['h3030]=8'h00; mem['h3031]=8'h00; mem['h3032]=8'h00; mem['h3033]=8'h00;
    mem['h3034]=8'h00; mem['h3035]=8'h00; mem['h3036]=8'h00; mem['h3037]=8'h00;
    mem['h3038]=8'h00; mem['h3039]=8'h00; mem['h303A]=8'h00; mem['h303B]=8'h00;
    mem['h303C]=8'h00; mem['h303D]=8'h00; mem['h303E]=8'h00; mem['h303F]=8'h00;
    mem['h3040]=8'h00; mem['h3041]=8'h00; mem['h3042]=8'h00; mem['h3043]=8'h00;
    mem['h3044]=8'h00; mem['h3045]=8'h00; mem['h3046]=8'h00; mem['h3047]=8'h00;
    mem['h3048]=8'h00; mem['h3049]=8'h00; mem['h304A]=8'h00; mem['h304B]=8'h00;
    mem['h304C]=8'h00; mem['h304D]=8'h00; mem['h304E]=8'h00; mem['h304F]=8'h00;
    mem['h3050]=8'h00; mem['h3051]=8'h00; mem['h3052]=8'h00; mem['h3053]=8'h00;
    mem['h3054]=8'h00; mem['h3055]=8'h00; mem['h3056]=8'h00; mem['h3057]=8'h00;
    mem['h3058]=8'h00; mem['h3059]=8'h00; mem['h305A]=8'h00; mem['h305B]=8'h00;
    mem['h305C]=8'h00; mem['h305D]=8'h00; mem['h305E]=8'h00; mem['h305F]=8'h00;
    mem['h3060]=8'h00; mem['h3061]=8'h00; mem['h3062]=8'h00; mem['h3063]=8'h00;
    mem['h3064]=8'h00; mem['h3065]=8'h00; mem['h3066]=8'h00; mem['h3067]=8'h00;
    mem['h3068]=8'h00; mem['h3069]=8'h00; mem['h306A]=8'h00; mem['h306B]=8'h00;
    mem['h306C]=8'h00; mem['h306D]=8'h00; mem['h306E]=8'h00; mem['h306F]=8'h00;
    mem['h3070]=8'h00; mem['h3071]=8'h00; mem['h3072]=8'h00; mem['h3073]=8'h00;
    mem['h3074]=8'h00; mem['h3075]=8'h00; mem['h3076]=8'h00; mem['h3077]=8'h00;
    mem['h3078]=8'h00; mem['h3079]=8'h00; mem['h307A]=8'h00; mem['h307B]=8'h00;
    mem['h307C]=8'h00; mem['h307D]=8'h00; mem['h307E]=8'h00; mem['h307F]=8'h00;
    mem['h3080]=8'h00; mem['h3081]=8'h00; mem['h3082]=8'h00; mem['h3083]=8'h00;
    mem['h3084]=8'h00; mem['h3085]=8'h00; mem['h3086]=8'h00; mem['h3087]=8'h00;
    mem['h3088]=8'h00; mem['h3089]=8'h00; mem['h308A]=8'h00; mem['h308B]=8'h00;
    mem['h308C]=8'h00; mem['h308D]=8'h00; mem['h308E]=8'h00; mem['h308F]=8'h00;
    mem['h3090]=8'h00; mem['h3091]=8'h00; mem['h3092]=8'h00; mem['h3093]=8'h00;
    mem['h3094]=8'h00; mem['h3095]=8'h00; mem['h3096]=8'h00; mem['h3097]=8'h00;
    mem['h3098]=8'h00; mem['h3099]=8'h00; mem['h309A]=8'h00; mem['h309B]=8'h00;
    mem['h309C]=8'h00; mem['h309D]=8'h00; mem['h309E]=8'h00; mem['h309F]=8'h00;
    mem['h30A0]=8'h00; mem['h30A1]=8'h00; mem['h30A2]=8'h00; mem['h30A3]=8'h00;
    mem['h30A4]=8'h00; mem['h30A5]=8'h00; mem['h30A6]=8'h00; mem['h30A7]=8'h00;
    mem['h30A8]=8'h00; mem['h30A9]=8'h00; mem['h30AA]=8'h00; mem['h30AB]=8'h00;
    mem['h30AC]=8'h00; mem['h30AD]=8'h00; mem['h30AE]=8'h00; mem['h30AF]=8'h00;
    mem['h30B0]=8'h00; mem['h30B1]=8'h00; mem['h30B2]=8'h00; mem['h30B3]=8'h00;
    mem['h30B4]=8'h00; mem['h30B5]=8'h00; mem['h30B6]=8'h00; mem['h30B7]=8'h00;
    mem['h30B8]=8'h00; mem['h30B9]=8'h00; mem['h30BA]=8'h00; mem['h30BB]=8'h00;
    mem['h30BC]=8'h00; mem['h30BD]=8'h00; mem['h30BE]=8'h00; mem['h30BF]=8'h00;
    mem['h30C0]=8'h00; mem['h30C1]=8'h00; mem['h30C2]=8'h00; mem['h30C3]=8'h00;
    mem['h30C4]=8'h00; mem['h30C5]=8'h00; mem['h30C6]=8'h00; mem['h30C7]=8'h00;
    mem['h30C8]=8'h00; mem['h30C9]=8'h00; mem['h30CA]=8'h00; mem['h30CB]=8'h00;
    mem['h30CC]=8'h00; mem['h30CD]=8'h00; mem['h30CE]=8'h00; mem['h30CF]=8'h00;
    mem['h30D0]=8'h00; mem['h30D1]=8'h00; mem['h30D2]=8'h00; mem['h30D3]=8'h00;
    mem['h30D4]=8'h00; mem['h30D5]=8'h00; mem['h30D6]=8'h00; mem['h30D7]=8'h00;
    mem['h30D8]=8'h00; mem['h30D9]=8'h00; mem['h30DA]=8'h00; mem['h30DB]=8'h00;
    mem['h30DC]=8'h00; mem['h30DD]=8'h00; mem['h30DE]=8'h00; mem['h30DF]=8'h00;
    mem['h30E0]=8'h00; mem['h30E1]=8'h00; mem['h30E2]=8'h00; mem['h30E3]=8'h00;
    mem['h30E4]=8'h00; mem['h30E5]=8'h00; mem['h30E6]=8'h00; mem['h30E7]=8'h00;
    mem['h30E8]=8'h00; mem['h30E9]=8'h00; mem['h30EA]=8'h00; mem['h30EB]=8'h00;
    mem['h30EC]=8'h00; mem['h30ED]=8'h00; mem['h30EE]=8'h00; mem['h30EF]=8'h00;
    mem['h30F0]=8'h00; mem['h30F1]=8'h00; mem['h30F2]=8'h00; mem['h30F3]=8'h00;
    mem['h30F4]=8'h00; mem['h30F5]=8'h00; mem['h30F6]=8'h00; mem['h30F7]=8'h00;
    mem['h30F8]=8'h00; mem['h30F9]=8'h00; mem['h30FA]=8'h00; mem['h30FB]=8'h00;
    mem['h30FC]=8'h00; mem['h30FD]=8'h00; mem['h30FE]=8'h00; mem['h30FF]=8'h00;
    mem['h3100]=8'h00; mem['h3101]=8'h00; mem['h3102]=8'h00; mem['h3103]=8'h00;
    mem['h3104]=8'h00; mem['h3105]=8'h00; mem['h3106]=8'h00; mem['h3107]=8'h00;
    mem['h3108]=8'h00; mem['h3109]=8'h00; mem['h310A]=8'h00; mem['h310B]=8'h00;
    mem['h310C]=8'h00; mem['h310D]=8'h00; mem['h310E]=8'h00; mem['h310F]=8'h00;
    mem['h3110]=8'h00; mem['h3111]=8'h00; mem['h3112]=8'h00; mem['h3113]=8'h00;
    mem['h3114]=8'h00; mem['h3115]=8'h00; mem['h3116]=8'h00; mem['h3117]=8'h00;
    mem['h3118]=8'h00; mem['h3119]=8'h00; mem['h311A]=8'h00; mem['h311B]=8'h00;
    mem['h311C]=8'h00; mem['h311D]=8'h00; mem['h311E]=8'h00; mem['h311F]=8'h00;
    mem['h3120]=8'h00; mem['h3121]=8'h00; mem['h3122]=8'h00; mem['h3123]=8'h00;
    mem['h3124]=8'h00; mem['h3125]=8'h00; mem['h3126]=8'h00; mem['h3127]=8'h00;
    mem['h3128]=8'h00; mem['h3129]=8'h00; mem['h312A]=8'h00; mem['h312B]=8'h00;
    mem['h312C]=8'h00; mem['h312D]=8'h00; mem['h312E]=8'h00; mem['h312F]=8'h00;
    mem['h3130]=8'h00; mem['h3131]=8'h00; mem['h3132]=8'h00; mem['h3133]=8'h00;
    mem['h3134]=8'h00; mem['h3135]=8'h00; mem['h3136]=8'h00; mem['h3137]=8'h00;
    mem['h3138]=8'h00; mem['h3139]=8'h00; mem['h313A]=8'h00; mem['h313B]=8'h00;
    mem['h313C]=8'h00; mem['h313D]=8'h00; mem['h313E]=8'h00; mem['h313F]=8'h00;
    mem['h3140]=8'h00; mem['h3141]=8'h00; mem['h3142]=8'h00; mem['h3143]=8'h00;
    mem['h3144]=8'h00; mem['h3145]=8'h00; mem['h3146]=8'h00; mem['h3147]=8'h00;
    mem['h3148]=8'h00; mem['h3149]=8'h00; mem['h314A]=8'h00; mem['h314B]=8'h00;
    mem['h314C]=8'h00; mem['h314D]=8'h00; mem['h314E]=8'h00; mem['h314F]=8'h00;
    mem['h3150]=8'h00; mem['h3151]=8'h00; mem['h3152]=8'h00; mem['h3153]=8'h00;
    mem['h3154]=8'h00; mem['h3155]=8'h00; mem['h3156]=8'h00; mem['h3157]=8'h00;
    mem['h3158]=8'h00; mem['h3159]=8'h00; mem['h315A]=8'h00; mem['h315B]=8'h00;
    mem['h315C]=8'h00; mem['h315D]=8'h00; mem['h315E]=8'h00; mem['h315F]=8'h00;
    mem['h3160]=8'h00; mem['h3161]=8'h00; mem['h3162]=8'h00; mem['h3163]=8'h00;
    mem['h3164]=8'h00; mem['h3165]=8'h00; mem['h3166]=8'h00; mem['h3167]=8'h00;
    mem['h3168]=8'h00; mem['h3169]=8'h00; mem['h316A]=8'h00; mem['h316B]=8'h00;
    mem['h316C]=8'h00; mem['h316D]=8'h00; mem['h316E]=8'h00; mem['h316F]=8'h00;
    mem['h3170]=8'h00; mem['h3171]=8'h00; mem['h3172]=8'h00; mem['h3173]=8'h00;
    mem['h3174]=8'h00; mem['h3175]=8'h00; mem['h3176]=8'h00; mem['h3177]=8'h00;
    mem['h3178]=8'h00; mem['h3179]=8'h00; mem['h317A]=8'h00; mem['h317B]=8'h00;
    mem['h317C]=8'h00; mem['h317D]=8'h00; mem['h317E]=8'h00; mem['h317F]=8'h00;
    mem['h3180]=8'h00; mem['h3181]=8'h00; mem['h3182]=8'h00; mem['h3183]=8'h00;
    mem['h3184]=8'h00; mem['h3185]=8'h00; mem['h3186]=8'h00; mem['h3187]=8'h00;
    mem['h3188]=8'h00; mem['h3189]=8'h00; mem['h318A]=8'h00; mem['h318B]=8'h00;
    mem['h318C]=8'h00; mem['h318D]=8'h00; mem['h318E]=8'h00; mem['h318F]=8'h00;
    mem['h3190]=8'h00; mem['h3191]=8'h00; mem['h3192]=8'h00; mem['h3193]=8'h00;
    mem['h3194]=8'h00; mem['h3195]=8'h00; mem['h3196]=8'h00; mem['h3197]=8'h00;
    mem['h3198]=8'h00; mem['h3199]=8'h00; mem['h319A]=8'h00; mem['h319B]=8'h00;
    mem['h319C]=8'h00; mem['h319D]=8'h00; mem['h319E]=8'h00; mem['h319F]=8'h00;
    mem['h31A0]=8'h00; mem['h31A1]=8'h00; mem['h31A2]=8'h00; mem['h31A3]=8'h00;
    mem['h31A4]=8'h00; mem['h31A5]=8'h00; mem['h31A6]=8'h00; mem['h31A7]=8'h00;
    mem['h31A8]=8'h00; mem['h31A9]=8'h00; mem['h31AA]=8'h00; mem['h31AB]=8'h00;
    mem['h31AC]=8'h00; mem['h31AD]=8'h00; mem['h31AE]=8'h00; mem['h31AF]=8'h00;
    mem['h31B0]=8'h00; mem['h31B1]=8'h00; mem['h31B2]=8'h00; mem['h31B3]=8'h00;
    mem['h31B4]=8'h00; mem['h31B5]=8'h00; mem['h31B6]=8'h00; mem['h31B7]=8'h00;
    mem['h31B8]=8'h00; mem['h31B9]=8'h00; mem['h31BA]=8'h00; mem['h31BB]=8'h00;
    mem['h31BC]=8'h00; mem['h31BD]=8'h00; mem['h31BE]=8'h00; mem['h31BF]=8'h00;
    mem['h31C0]=8'h00; mem['h31C1]=8'h00; mem['h31C2]=8'h00; mem['h31C3]=8'h00;
    mem['h31C4]=8'h00; mem['h31C5]=8'h00; mem['h31C6]=8'h00; mem['h31C7]=8'h00;
    mem['h31C8]=8'h00; mem['h31C9]=8'h00; mem['h31CA]=8'h00; mem['h31CB]=8'h00;
    mem['h31CC]=8'h00; mem['h31CD]=8'h00; mem['h31CE]=8'h00; mem['h31CF]=8'h00;
    mem['h31D0]=8'h00; mem['h31D1]=8'h00; mem['h31D2]=8'h00; mem['h31D3]=8'h00;
    mem['h31D4]=8'h00; mem['h31D5]=8'h00; mem['h31D6]=8'h00; mem['h31D7]=8'h00;
    mem['h31D8]=8'h00; mem['h31D9]=8'h00; mem['h31DA]=8'h00; mem['h31DB]=8'h00;
    mem['h31DC]=8'h00; mem['h31DD]=8'h00; mem['h31DE]=8'h00; mem['h31DF]=8'h00;
    mem['h31E0]=8'h00; mem['h31E1]=8'h00; mem['h31E2]=8'h00; mem['h31E3]=8'h00;
    mem['h31E4]=8'h00; mem['h31E5]=8'h00; mem['h31E6]=8'h00; mem['h31E7]=8'h00;
    mem['h31E8]=8'h00; mem['h31E9]=8'h00; mem['h31EA]=8'h00; mem['h31EB]=8'h00;
    mem['h31EC]=8'h00; mem['h31ED]=8'h00; mem['h31EE]=8'h00; mem['h31EF]=8'h00;
    mem['h31F0]=8'h00; mem['h31F1]=8'h00; mem['h31F2]=8'h00; mem['h31F3]=8'h00;
    mem['h31F4]=8'h00; mem['h31F5]=8'h00; mem['h31F6]=8'h00; mem['h31F7]=8'h00;
    mem['h31F8]=8'h00; mem['h31F9]=8'h00; mem['h31FA]=8'h00; mem['h31FB]=8'h00;
    mem['h31FC]=8'h00; mem['h31FD]=8'h00; mem['h31FE]=8'h00; mem['h31FF]=8'h00;
    mem['h3200]=8'h00; mem['h3201]=8'h00; mem['h3202]=8'h00; mem['h3203]=8'h00;
    mem['h3204]=8'h00; mem['h3205]=8'h00; mem['h3206]=8'h00; mem['h3207]=8'h00;
    mem['h3208]=8'h00; mem['h3209]=8'h00; mem['h320A]=8'h00; mem['h320B]=8'h00;
    mem['h320C]=8'h00; mem['h320D]=8'h00; mem['h320E]=8'h00; mem['h320F]=8'h00;
    mem['h3210]=8'h00; mem['h3211]=8'h00; mem['h3212]=8'h00; mem['h3213]=8'h00;
    mem['h3214]=8'h00; mem['h3215]=8'h00; mem['h3216]=8'h00; mem['h3217]=8'h00;
    mem['h3218]=8'h00; mem['h3219]=8'h00; mem['h321A]=8'h00; mem['h321B]=8'h00;
    mem['h321C]=8'h00; mem['h321D]=8'h00; mem['h321E]=8'h00; mem['h321F]=8'h00;
    mem['h3220]=8'h00; mem['h3221]=8'h00; mem['h3222]=8'h00; mem['h3223]=8'h00;
    mem['h3224]=8'h00; mem['h3225]=8'h00; mem['h3226]=8'h00; mem['h3227]=8'h00;
    mem['h3228]=8'h00; mem['h3229]=8'h00; mem['h322A]=8'h00; mem['h322B]=8'h00;
    mem['h322C]=8'h00; mem['h322D]=8'h00; mem['h322E]=8'h00; mem['h322F]=8'h00;
    mem['h3230]=8'h00; mem['h3231]=8'h00; mem['h3232]=8'h00; mem['h3233]=8'h00;
    mem['h3234]=8'h00; mem['h3235]=8'h00; mem['h3236]=8'h00; mem['h3237]=8'h00;
    mem['h3238]=8'h00; mem['h3239]=8'h00; mem['h323A]=8'h00; mem['h323B]=8'h00;
    mem['h323C]=8'h00; mem['h323D]=8'h00; mem['h323E]=8'h00; mem['h323F]=8'h00;
    mem['h3240]=8'h00; mem['h3241]=8'h00; mem['h3242]=8'h00; mem['h3243]=8'h00;
    mem['h3244]=8'h00; mem['h3245]=8'h00; mem['h3246]=8'h00; mem['h3247]=8'h00;
    mem['h3248]=8'h00; mem['h3249]=8'h00; mem['h324A]=8'h00; mem['h324B]=8'h00;
    mem['h324C]=8'h00; mem['h324D]=8'h00; mem['h324E]=8'h00; mem['h324F]=8'h00;
    mem['h3250]=8'h00; mem['h3251]=8'h00; mem['h3252]=8'h00; mem['h3253]=8'h00;
    mem['h3254]=8'h00; mem['h3255]=8'h00; mem['h3256]=8'h00; mem['h3257]=8'h00;
    mem['h3258]=8'h00; mem['h3259]=8'h00; mem['h325A]=8'h00; mem['h325B]=8'h00;
    mem['h325C]=8'h00; mem['h325D]=8'h00; mem['h325E]=8'h00; mem['h325F]=8'h00;
    mem['h3260]=8'h00; mem['h3261]=8'h00; mem['h3262]=8'h00; mem['h3263]=8'h00;
    mem['h3264]=8'h00; mem['h3265]=8'h00; mem['h3266]=8'h00; mem['h3267]=8'h00;
    mem['h3268]=8'h00; mem['h3269]=8'h00; mem['h326A]=8'h00; mem['h326B]=8'h00;
    mem['h326C]=8'h00; mem['h326D]=8'h00; mem['h326E]=8'h00; mem['h326F]=8'h00;
    mem['h3270]=8'h00; mem['h3271]=8'h00; mem['h3272]=8'h00; mem['h3273]=8'h00;
    mem['h3274]=8'h00; mem['h3275]=8'h00; mem['h3276]=8'h00; mem['h3277]=8'h00;
    mem['h3278]=8'h00; mem['h3279]=8'h00; mem['h327A]=8'h00; mem['h327B]=8'h00;
    mem['h327C]=8'h00; mem['h327D]=8'h00; mem['h327E]=8'h00; mem['h327F]=8'h00;
    mem['h3280]=8'h00; mem['h3281]=8'h00; mem['h3282]=8'h00; mem['h3283]=8'h00;
    mem['h3284]=8'h00; mem['h3285]=8'h00; mem['h3286]=8'h00; mem['h3287]=8'h00;
    mem['h3288]=8'h00; mem['h3289]=8'h00; mem['h328A]=8'h00; mem['h328B]=8'h00;
    mem['h328C]=8'h00; mem['h328D]=8'h00; mem['h328E]=8'h00; mem['h328F]=8'h00;
    mem['h3290]=8'h00; mem['h3291]=8'h00; mem['h3292]=8'h00; mem['h3293]=8'h00;
    mem['h3294]=8'h00; mem['h3295]=8'h00; mem['h3296]=8'h00; mem['h3297]=8'h00;
    mem['h3298]=8'h00; mem['h3299]=8'h00; mem['h329A]=8'h00; mem['h329B]=8'h00;
    mem['h329C]=8'h00; mem['h329D]=8'h00; mem['h329E]=8'h00; mem['h329F]=8'h00;
    mem['h32A0]=8'h00; mem['h32A1]=8'h00; mem['h32A2]=8'h00; mem['h32A3]=8'h00;
    mem['h32A4]=8'h00; mem['h32A5]=8'h00; mem['h32A6]=8'h00; mem['h32A7]=8'h00;
    mem['h32A8]=8'h00; mem['h32A9]=8'h00; mem['h32AA]=8'h00; mem['h32AB]=8'h00;
    mem['h32AC]=8'h00; mem['h32AD]=8'h00; mem['h32AE]=8'h00; mem['h32AF]=8'h00;
    mem['h32B0]=8'h00; mem['h32B1]=8'h00; mem['h32B2]=8'h00; mem['h32B3]=8'h00;
    mem['h32B4]=8'h00; mem['h32B5]=8'h00; mem['h32B6]=8'h00; mem['h32B7]=8'h00;
    mem['h32B8]=8'h00; mem['h32B9]=8'h00; mem['h32BA]=8'h00; mem['h32BB]=8'h00;
    mem['h32BC]=8'h00; mem['h32BD]=8'h00; mem['h32BE]=8'h00; mem['h32BF]=8'h00;
    mem['h32C0]=8'h00; mem['h32C1]=8'h00; mem['h32C2]=8'h00; mem['h32C3]=8'h00;
    mem['h32C4]=8'h00; mem['h32C5]=8'h00; mem['h32C6]=8'h00; mem['h32C7]=8'h00;
    mem['h32C8]=8'h00; mem['h32C9]=8'h00; mem['h32CA]=8'h00; mem['h32CB]=8'h00;
    mem['h32CC]=8'h00; mem['h32CD]=8'h00; mem['h32CE]=8'h00; mem['h32CF]=8'h00;
    mem['h32D0]=8'h00; mem['h32D1]=8'h00; mem['h32D2]=8'h00; mem['h32D3]=8'h00;
    mem['h32D4]=8'h00; mem['h32D5]=8'h00; mem['h32D6]=8'h00; mem['h32D7]=8'h00;
    mem['h32D8]=8'h00; mem['h32D9]=8'h00; mem['h32DA]=8'h00; mem['h32DB]=8'h00;
    mem['h32DC]=8'h00; mem['h32DD]=8'h00; mem['h32DE]=8'h00; mem['h32DF]=8'h00;
    mem['h32E0]=8'h00; mem['h32E1]=8'h00; mem['h32E2]=8'h00; mem['h32E3]=8'h00;
    mem['h32E4]=8'h00; mem['h32E5]=8'h00; mem['h32E6]=8'h00; mem['h32E7]=8'h00;
    mem['h32E8]=8'h00; mem['h32E9]=8'h00; mem['h32EA]=8'h00; mem['h32EB]=8'h00;
    mem['h32EC]=8'h00; mem['h32ED]=8'h00; mem['h32EE]=8'h00; mem['h32EF]=8'h00;
    mem['h32F0]=8'h00; mem['h32F1]=8'h00; mem['h32F2]=8'h00; mem['h32F3]=8'h00;
    mem['h32F4]=8'h00; mem['h32F5]=8'h00; mem['h32F6]=8'h00; mem['h32F7]=8'h00;
    mem['h32F8]=8'h00; mem['h32F9]=8'h00; mem['h32FA]=8'h00; mem['h32FB]=8'h00;
    mem['h32FC]=8'h00; mem['h32FD]=8'h00; mem['h32FE]=8'h00; mem['h32FF]=8'h00;
    mem['h3300]=8'h00; mem['h3301]=8'h00; mem['h3302]=8'h00; mem['h3303]=8'h00;
    mem['h3304]=8'h00; mem['h3305]=8'h00; mem['h3306]=8'h00; mem['h3307]=8'h00;
    mem['h3308]=8'h00; mem['h3309]=8'h00; mem['h330A]=8'h00; mem['h330B]=8'h00;
    mem['h330C]=8'h00; mem['h330D]=8'h00; mem['h330E]=8'h00; mem['h330F]=8'h00;
    mem['h3310]=8'h00; mem['h3311]=8'h00; mem['h3312]=8'h00; mem['h3313]=8'h00;
    mem['h3314]=8'h00; mem['h3315]=8'h00; mem['h3316]=8'h00; mem['h3317]=8'h00;
    mem['h3318]=8'h00; mem['h3319]=8'h00; mem['h331A]=8'h00; mem['h331B]=8'h00;
    mem['h331C]=8'h00; mem['h331D]=8'h00; mem['h331E]=8'h00; mem['h331F]=8'h00;
    mem['h3320]=8'h00; mem['h3321]=8'h00; mem['h3322]=8'h00; mem['h3323]=8'h00;
    mem['h3324]=8'h00; mem['h3325]=8'h00; mem['h3326]=8'h00; mem['h3327]=8'h00;
    mem['h3328]=8'h00; mem['h3329]=8'h00; mem['h332A]=8'h00; mem['h332B]=8'h00;
    mem['h332C]=8'h00; mem['h332D]=8'h00; mem['h332E]=8'h00; mem['h332F]=8'h00;
    mem['h3330]=8'h00; mem['h3331]=8'h00; mem['h3332]=8'h00; mem['h3333]=8'h00;
    mem['h3334]=8'h00; mem['h3335]=8'h00; mem['h3336]=8'h00; mem['h3337]=8'h00;
    mem['h3338]=8'h00; mem['h3339]=8'h00; mem['h333A]=8'h00; mem['h333B]=8'h00;
    mem['h333C]=8'h00; mem['h333D]=8'h00; mem['h333E]=8'h00; mem['h333F]=8'h00;
    mem['h3340]=8'h00; mem['h3341]=8'h00; mem['h3342]=8'h00; mem['h3343]=8'h00;
    mem['h3344]=8'h00; mem['h3345]=8'h00; mem['h3346]=8'h00; mem['h3347]=8'h00;
    mem['h3348]=8'h00; mem['h3349]=8'h00; mem['h334A]=8'h00; mem['h334B]=8'h00;
    mem['h334C]=8'h00; mem['h334D]=8'h00; mem['h334E]=8'h00; mem['h334F]=8'h00;
    mem['h3350]=8'h00; mem['h3351]=8'h00; mem['h3352]=8'h00; mem['h3353]=8'h00;
    mem['h3354]=8'h00; mem['h3355]=8'h00; mem['h3356]=8'h00; mem['h3357]=8'h00;
    mem['h3358]=8'h00; mem['h3359]=8'h00; mem['h335A]=8'h00; mem['h335B]=8'h00;
    mem['h335C]=8'h00; mem['h335D]=8'h00; mem['h335E]=8'h00; mem['h335F]=8'h00;
    mem['h3360]=8'h00; mem['h3361]=8'h00; mem['h3362]=8'h00; mem['h3363]=8'h00;
    mem['h3364]=8'h00; mem['h3365]=8'h00; mem['h3366]=8'h00; mem['h3367]=8'h00;
    mem['h3368]=8'h00; mem['h3369]=8'h00; mem['h336A]=8'h00; mem['h336B]=8'h00;
    mem['h336C]=8'h00; mem['h336D]=8'h00; mem['h336E]=8'h00; mem['h336F]=8'h00;
    mem['h3370]=8'h00; mem['h3371]=8'h00; mem['h3372]=8'h00; mem['h3373]=8'h00;
    mem['h3374]=8'h00; mem['h3375]=8'h00; mem['h3376]=8'h00; mem['h3377]=8'h00;
    mem['h3378]=8'h00; mem['h3379]=8'h00; mem['h337A]=8'h00; mem['h337B]=8'h00;
    mem['h337C]=8'h00; mem['h337D]=8'h00; mem['h337E]=8'h00; mem['h337F]=8'h00;
    mem['h3380]=8'h00; mem['h3381]=8'h00; mem['h3382]=8'h00; mem['h3383]=8'h00;
    mem['h3384]=8'h00; mem['h3385]=8'h00; mem['h3386]=8'h00; mem['h3387]=8'h00;
    mem['h3388]=8'h00; mem['h3389]=8'h00; mem['h338A]=8'h00; mem['h338B]=8'h00;
    mem['h338C]=8'h00; mem['h338D]=8'h00; mem['h338E]=8'h00; mem['h338F]=8'h00;
    mem['h3390]=8'h00; mem['h3391]=8'h00; mem['h3392]=8'h00; mem['h3393]=8'h00;
    mem['h3394]=8'h00; mem['h3395]=8'h00; mem['h3396]=8'h00; mem['h3397]=8'h00;
    mem['h3398]=8'h00; mem['h3399]=8'h00; mem['h339A]=8'h00; mem['h339B]=8'h00;
    mem['h339C]=8'h00; mem['h339D]=8'h00; mem['h339E]=8'h00; mem['h339F]=8'h00;
    mem['h33A0]=8'h00; mem['h33A1]=8'h00; mem['h33A2]=8'h00; mem['h33A3]=8'h00;
    mem['h33A4]=8'h00; mem['h33A5]=8'h00; mem['h33A6]=8'h00; mem['h33A7]=8'h00;
    mem['h33A8]=8'h00; mem['h33A9]=8'h00; mem['h33AA]=8'h00; mem['h33AB]=8'h00;
    mem['h33AC]=8'h00; mem['h33AD]=8'h00; mem['h33AE]=8'h00; mem['h33AF]=8'h00;
    mem['h33B0]=8'h00; mem['h33B1]=8'h00; mem['h33B2]=8'h00; mem['h33B3]=8'h00;
    mem['h33B4]=8'h00; mem['h33B5]=8'h00; mem['h33B6]=8'h00; mem['h33B7]=8'h00;
    mem['h33B8]=8'h00; mem['h33B9]=8'h00; mem['h33BA]=8'h00; mem['h33BB]=8'h00;
    mem['h33BC]=8'h00; mem['h33BD]=8'h00; mem['h33BE]=8'h00; mem['h33BF]=8'h00;
    mem['h33C0]=8'h00; mem['h33C1]=8'h00; mem['h33C2]=8'h00; mem['h33C3]=8'h00;
    mem['h33C4]=8'h00; mem['h33C5]=8'h00; mem['h33C6]=8'h00; mem['h33C7]=8'h00;
    mem['h33C8]=8'h00; mem['h33C9]=8'h00; mem['h33CA]=8'h00; mem['h33CB]=8'h00;
    mem['h33CC]=8'h00; mem['h33CD]=8'h00; mem['h33CE]=8'h00; mem['h33CF]=8'h00;
    mem['h33D0]=8'h00; mem['h33D1]=8'h00; mem['h33D2]=8'h00; mem['h33D3]=8'h00;
    mem['h33D4]=8'h00; mem['h33D5]=8'h00; mem['h33D6]=8'h00; mem['h33D7]=8'h00;
    mem['h33D8]=8'h00; mem['h33D9]=8'h00; mem['h33DA]=8'h00; mem['h33DB]=8'h00;
    mem['h33DC]=8'h00; mem['h33DD]=8'h00; mem['h33DE]=8'h00; mem['h33DF]=8'h00;
    mem['h33E0]=8'h00; mem['h33E1]=8'h00; mem['h33E2]=8'h00; mem['h33E3]=8'h00;
    mem['h33E4]=8'h00; mem['h33E5]=8'h00; mem['h33E6]=8'h00; mem['h33E7]=8'h00;
    mem['h33E8]=8'h00; mem['h33E9]=8'h00; mem['h33EA]=8'h00; mem['h33EB]=8'h00;
    mem['h33EC]=8'h00; mem['h33ED]=8'h00; mem['h33EE]=8'h00; mem['h33EF]=8'h00;
    mem['h33F0]=8'h00; mem['h33F1]=8'h00; mem['h33F2]=8'h00; mem['h33F3]=8'h00;
    mem['h33F4]=8'h00; mem['h33F5]=8'h00; mem['h33F6]=8'h00; mem['h33F7]=8'h00;
    mem['h33F8]=8'h00; mem['h33F9]=8'h00; mem['h33FA]=8'h00; mem['h33FB]=8'h00;
    mem['h33FC]=8'h00; mem['h33FD]=8'h00; mem['h33FE]=8'h00; mem['h33FF]=8'h00;
    mem['h3400]=8'h00; mem['h3401]=8'h00; mem['h3402]=8'h00; mem['h3403]=8'h00;
    mem['h3404]=8'h00; mem['h3405]=8'h00; mem['h3406]=8'h00; mem['h3407]=8'h00;
    mem['h3408]=8'h00; mem['h3409]=8'h00; mem['h340A]=8'h00; mem['h340B]=8'h00;
    mem['h340C]=8'h00; mem['h340D]=8'h00; mem['h340E]=8'h00; mem['h340F]=8'h00;
    mem['h3410]=8'h00; mem['h3411]=8'h00; mem['h3412]=8'h00; mem['h3413]=8'h00;
    mem['h3414]=8'h00; mem['h3415]=8'h00; mem['h3416]=8'h00; mem['h3417]=8'h00;
    mem['h3418]=8'h00; mem['h3419]=8'h00; mem['h341A]=8'h00; mem['h341B]=8'h00;
    mem['h341C]=8'h00; mem['h341D]=8'h00; mem['h341E]=8'h00; mem['h341F]=8'h00;
    mem['h3420]=8'h00; mem['h3421]=8'h00; mem['h3422]=8'h00; mem['h3423]=8'h00;
    mem['h3424]=8'h00; mem['h3425]=8'h00; mem['h3426]=8'h00; mem['h3427]=8'h00;
    mem['h3428]=8'h00; mem['h3429]=8'h00; mem['h342A]=8'h00; mem['h342B]=8'h00;
    mem['h342C]=8'h00; mem['h342D]=8'h00; mem['h342E]=8'h00; mem['h342F]=8'h00;
    mem['h3430]=8'h00; mem['h3431]=8'h00; mem['h3432]=8'h00; mem['h3433]=8'h00;
    mem['h3434]=8'h00; mem['h3435]=8'h00; mem['h3436]=8'h00; mem['h3437]=8'h00;
    mem['h3438]=8'h00; mem['h3439]=8'h00; mem['h343A]=8'h00; mem['h343B]=8'h00;
    mem['h343C]=8'h00; mem['h343D]=8'h00; mem['h343E]=8'h00; mem['h343F]=8'h00;
    mem['h3440]=8'h00; mem['h3441]=8'h00; mem['h3442]=8'h00; mem['h3443]=8'h00;
    mem['h3444]=8'h00; mem['h3445]=8'h00; mem['h3446]=8'h00; mem['h3447]=8'h00;
    mem['h3448]=8'h00; mem['h3449]=8'h00; mem['h344A]=8'h00; mem['h344B]=8'h00;
    mem['h344C]=8'h00; mem['h344D]=8'h00; mem['h344E]=8'h00; mem['h344F]=8'h00;
    mem['h3450]=8'h00; mem['h3451]=8'h00; mem['h3452]=8'h00; mem['h3453]=8'h00;
    mem['h3454]=8'h00; mem['h3455]=8'h00; mem['h3456]=8'h00; mem['h3457]=8'h00;
    mem['h3458]=8'h00; mem['h3459]=8'h00; mem['h345A]=8'h00; mem['h345B]=8'h00;
    mem['h345C]=8'h00; mem['h345D]=8'h00; mem['h345E]=8'h00; mem['h345F]=8'h00;
    mem['h3460]=8'h00; mem['h3461]=8'h00; mem['h3462]=8'h00; mem['h3463]=8'h00;
    mem['h3464]=8'h00; mem['h3465]=8'h00; mem['h3466]=8'h00; mem['h3467]=8'h00;
    mem['h3468]=8'h00; mem['h3469]=8'h00; mem['h346A]=8'h00; mem['h346B]=8'h00;
    mem['h346C]=8'h00; mem['h346D]=8'h00; mem['h346E]=8'h00; mem['h346F]=8'h00;
    mem['h3470]=8'h00; mem['h3471]=8'h00; mem['h3472]=8'h00; mem['h3473]=8'h00;
    mem['h3474]=8'h00; mem['h3475]=8'h00; mem['h3476]=8'h00; mem['h3477]=8'h00;
    mem['h3478]=8'h00; mem['h3479]=8'h00; mem['h347A]=8'h00; mem['h347B]=8'h00;
    mem['h347C]=8'h00; mem['h347D]=8'h00; mem['h347E]=8'h00; mem['h347F]=8'h00;
    mem['h3480]=8'h00; mem['h3481]=8'h00; mem['h3482]=8'h00; mem['h3483]=8'h00;
    mem['h3484]=8'h00; mem['h3485]=8'h00; mem['h3486]=8'h00; mem['h3487]=8'h00;
    mem['h3488]=8'h00; mem['h3489]=8'h00; mem['h348A]=8'h00; mem['h348B]=8'h00;
    mem['h348C]=8'h00; mem['h348D]=8'h00; mem['h348E]=8'h00; mem['h348F]=8'h00;
    mem['h3490]=8'h00; mem['h3491]=8'h00; mem['h3492]=8'h00; mem['h3493]=8'h00;
    mem['h3494]=8'h00; mem['h3495]=8'h00; mem['h3496]=8'h00; mem['h3497]=8'h00;
    mem['h3498]=8'h00; mem['h3499]=8'h00; mem['h349A]=8'h00; mem['h349B]=8'h00;
    mem['h349C]=8'h00; mem['h349D]=8'h00; mem['h349E]=8'h00; mem['h349F]=8'h00;
    mem['h34A0]=8'h00; mem['h34A1]=8'h00; mem['h34A2]=8'h00; mem['h34A3]=8'h00;
    mem['h34A4]=8'h00; mem['h34A5]=8'h00; mem['h34A6]=8'h00; mem['h34A7]=8'h00;
    mem['h34A8]=8'h00; mem['h34A9]=8'h00; mem['h34AA]=8'h00; mem['h34AB]=8'h00;
    mem['h34AC]=8'h00; mem['h34AD]=8'h00; mem['h34AE]=8'h00; mem['h34AF]=8'h00;
    mem['h34B0]=8'h00; mem['h34B1]=8'h00; mem['h34B2]=8'h00; mem['h34B3]=8'h00;
    mem['h34B4]=8'h00; mem['h34B5]=8'h00; mem['h34B6]=8'h00; mem['h34B7]=8'h00;
    mem['h34B8]=8'h00; mem['h34B9]=8'h00; mem['h34BA]=8'h00; mem['h34BB]=8'h00;
    mem['h34BC]=8'h00; mem['h34BD]=8'h00; mem['h34BE]=8'h00; mem['h34BF]=8'h00;
    mem['h34C0]=8'h00; mem['h34C1]=8'h00; mem['h34C2]=8'h00; mem['h34C3]=8'h00;
    mem['h34C4]=8'h00; mem['h34C5]=8'h00; mem['h34C6]=8'h00; mem['h34C7]=8'h00;
    mem['h34C8]=8'h00; mem['h34C9]=8'h00; mem['h34CA]=8'h00; mem['h34CB]=8'h00;
    mem['h34CC]=8'h00; mem['h34CD]=8'h00; mem['h34CE]=8'h00; mem['h34CF]=8'h00;
    mem['h34D0]=8'h00; mem['h34D1]=8'h00; mem['h34D2]=8'h00; mem['h34D3]=8'h00;
    mem['h34D4]=8'h00; mem['h34D5]=8'h00; mem['h34D6]=8'h00; mem['h34D7]=8'h00;
    mem['h34D8]=8'h00; mem['h34D9]=8'h00; mem['h34DA]=8'h00; mem['h34DB]=8'h00;
    mem['h34DC]=8'h00; mem['h34DD]=8'h00; mem['h34DE]=8'h00; mem['h34DF]=8'h00;
    mem['h34E0]=8'h00; mem['h34E1]=8'h00; mem['h34E2]=8'h00; mem['h34E3]=8'h00;
    mem['h34E4]=8'h00; mem['h34E5]=8'h00; mem['h34E6]=8'h00; mem['h34E7]=8'h00;
    mem['h34E8]=8'h00; mem['h34E9]=8'h00; mem['h34EA]=8'h00; mem['h34EB]=8'h00;
    mem['h34EC]=8'h00; mem['h34ED]=8'h00; mem['h34EE]=8'h00; mem['h34EF]=8'h00;
    mem['h34F0]=8'h00; mem['h34F1]=8'h00; mem['h34F2]=8'h00; mem['h34F3]=8'h00;
    mem['h34F4]=8'h00; mem['h34F5]=8'h00; mem['h34F6]=8'h00; mem['h34F7]=8'h00;
    mem['h34F8]=8'h00; mem['h34F9]=8'h00; mem['h34FA]=8'h00; mem['h34FB]=8'h00;
    mem['h34FC]=8'h00; mem['h34FD]=8'h00; mem['h34FE]=8'h00; mem['h34FF]=8'h00;
    mem['h3500]=8'h00; mem['h3501]=8'h00; mem['h3502]=8'h00; mem['h3503]=8'h00;
    mem['h3504]=8'h00; mem['h3505]=8'h00; mem['h3506]=8'h00; mem['h3507]=8'h00;
    mem['h3508]=8'h00; mem['h3509]=8'h00; mem['h350A]=8'h00; mem['h350B]=8'h00;
    mem['h350C]=8'h00; mem['h350D]=8'h00; mem['h350E]=8'h00; mem['h350F]=8'h00;
    mem['h3510]=8'h00; mem['h3511]=8'h00; mem['h3512]=8'h00; mem['h3513]=8'h00;
    mem['h3514]=8'h00; mem['h3515]=8'h00; mem['h3516]=8'h00; mem['h3517]=8'h00;
    mem['h3518]=8'h00; mem['h3519]=8'h00; mem['h351A]=8'h00; mem['h351B]=8'h00;
    mem['h351C]=8'h00; mem['h351D]=8'h00; mem['h351E]=8'h00; mem['h351F]=8'h00;
    mem['h3520]=8'h00; mem['h3521]=8'h00; mem['h3522]=8'h00; mem['h3523]=8'h00;
    mem['h3524]=8'h00; mem['h3525]=8'h00; mem['h3526]=8'h00; mem['h3527]=8'h00;
    mem['h3528]=8'h00; mem['h3529]=8'h00; mem['h352A]=8'h00; mem['h352B]=8'h00;
    mem['h352C]=8'h00; mem['h352D]=8'h00; mem['h352E]=8'h00; mem['h352F]=8'h00;
    mem['h3530]=8'h00; mem['h3531]=8'h00; mem['h3532]=8'h00; mem['h3533]=8'h00;
    mem['h3534]=8'h00; mem['h3535]=8'h00; mem['h3536]=8'h00; mem['h3537]=8'h00;
    mem['h3538]=8'h00; mem['h3539]=8'h00; mem['h353A]=8'h00; mem['h353B]=8'h00;
    mem['h353C]=8'h00; mem['h353D]=8'h00; mem['h353E]=8'h00; mem['h353F]=8'h00;
    mem['h3540]=8'h00; mem['h3541]=8'h00; mem['h3542]=8'h00; mem['h3543]=8'h00;
    mem['h3544]=8'h00; mem['h3545]=8'h00; mem['h3546]=8'h00; mem['h3547]=8'h00;
    mem['h3548]=8'h00; mem['h3549]=8'h00; mem['h354A]=8'h00; mem['h354B]=8'h00;
    mem['h354C]=8'h00; mem['h354D]=8'h00; mem['h354E]=8'h00; mem['h354F]=8'h00;
    mem['h3550]=8'h00; mem['h3551]=8'h00; mem['h3552]=8'h00; mem['h3553]=8'h00;
    mem['h3554]=8'h00; mem['h3555]=8'h00; mem['h3556]=8'h00; mem['h3557]=8'h00;
    mem['h3558]=8'h00; mem['h3559]=8'h00; mem['h355A]=8'h00; mem['h355B]=8'h00;
    mem['h355C]=8'h00; mem['h355D]=8'h00; mem['h355E]=8'h00; mem['h355F]=8'h00;
    mem['h3560]=8'h00; mem['h3561]=8'h00; mem['h3562]=8'h00; mem['h3563]=8'h00;
    mem['h3564]=8'h00; mem['h3565]=8'h00; mem['h3566]=8'h00; mem['h3567]=8'h00;
    mem['h3568]=8'h00; mem['h3569]=8'h00; mem['h356A]=8'h00; mem['h356B]=8'h00;
    mem['h356C]=8'h00; mem['h356D]=8'h00; mem['h356E]=8'h00; mem['h356F]=8'h00;
    mem['h3570]=8'h00; mem['h3571]=8'h00; mem['h3572]=8'h00; mem['h3573]=8'h00;
    mem['h3574]=8'h00; mem['h3575]=8'h00; mem['h3576]=8'h00; mem['h3577]=8'h00;
    mem['h3578]=8'h00; mem['h3579]=8'h00; mem['h357A]=8'h00; mem['h357B]=8'h00;
    mem['h357C]=8'h00; mem['h357D]=8'h00; mem['h357E]=8'h00; mem['h357F]=8'h00;
    mem['h3580]=8'h00; mem['h3581]=8'h00; mem['h3582]=8'h00; mem['h3583]=8'h00;
    mem['h3584]=8'h00; mem['h3585]=8'h00; mem['h3586]=8'h00; mem['h3587]=8'h00;
    mem['h3588]=8'h00; mem['h3589]=8'h00; mem['h358A]=8'h00; mem['h358B]=8'h00;
    mem['h358C]=8'h00; mem['h358D]=8'h00; mem['h358E]=8'h00; mem['h358F]=8'h00;
    mem['h3590]=8'h00; mem['h3591]=8'h00; mem['h3592]=8'h00; mem['h3593]=8'h00;
    mem['h3594]=8'h00; mem['h3595]=8'h00; mem['h3596]=8'h00; mem['h3597]=8'h00;
    mem['h3598]=8'h00; mem['h3599]=8'h00; mem['h359A]=8'h00; mem['h359B]=8'h00;
    mem['h359C]=8'h00; mem['h359D]=8'h00; mem['h359E]=8'h00; mem['h359F]=8'h00;
    mem['h35A0]=8'h00; mem['h35A1]=8'h00; mem['h35A2]=8'h00; mem['h35A3]=8'h00;
    mem['h35A4]=8'h00; mem['h35A5]=8'h00; mem['h35A6]=8'h00; mem['h35A7]=8'h00;
    mem['h35A8]=8'h00; mem['h35A9]=8'h00; mem['h35AA]=8'h00; mem['h35AB]=8'h00;
    mem['h35AC]=8'h00; mem['h35AD]=8'h00; mem['h35AE]=8'h00; mem['h35AF]=8'h00;
    mem['h35B0]=8'h00; mem['h35B1]=8'h00; mem['h35B2]=8'h00; mem['h35B3]=8'h00;
    mem['h35B4]=8'h00; mem['h35B5]=8'h00; mem['h35B6]=8'h00; mem['h35B7]=8'h00;
    mem['h35B8]=8'h00; mem['h35B9]=8'h00; mem['h35BA]=8'h00; mem['h35BB]=8'h00;
    mem['h35BC]=8'h00; mem['h35BD]=8'h00; mem['h35BE]=8'h00; mem['h35BF]=8'h00;
    mem['h35C0]=8'h00; mem['h35C1]=8'h00; mem['h35C2]=8'h00; mem['h35C3]=8'h00;
    mem['h35C4]=8'h00; mem['h35C5]=8'h00; mem['h35C6]=8'h00; mem['h35C7]=8'h00;
    mem['h35C8]=8'h00; mem['h35C9]=8'h00; mem['h35CA]=8'h00; mem['h35CB]=8'h00;
    mem['h35CC]=8'h00; mem['h35CD]=8'h00; mem['h35CE]=8'h00; mem['h35CF]=8'h00;
    mem['h35D0]=8'h00; mem['h35D1]=8'h00; mem['h35D2]=8'h00; mem['h35D3]=8'h00;
    mem['h35D4]=8'h00; mem['h35D5]=8'h00; mem['h35D6]=8'h00; mem['h35D7]=8'h00;
    mem['h35D8]=8'h00; mem['h35D9]=8'h00; mem['h35DA]=8'h00; mem['h35DB]=8'h00;
    mem['h35DC]=8'h00; mem['h35DD]=8'h00; mem['h35DE]=8'h00; mem['h35DF]=8'h00;
    mem['h35E0]=8'h00; mem['h35E1]=8'h00; mem['h35E2]=8'h00; mem['h35E3]=8'h00;
    mem['h35E4]=8'h00; mem['h35E5]=8'h00; mem['h35E6]=8'h00; mem['h35E7]=8'h00;
    mem['h35E8]=8'h00; mem['h35E9]=8'h00; mem['h35EA]=8'h00; mem['h35EB]=8'h00;
    mem['h35EC]=8'h00; mem['h35ED]=8'h00; mem['h35EE]=8'h00; mem['h35EF]=8'h00;
    mem['h35F0]=8'h00; mem['h35F1]=8'h00; mem['h35F2]=8'h00; mem['h35F3]=8'h00;
    mem['h35F4]=8'h00; mem['h35F5]=8'h00; mem['h35F6]=8'h00; mem['h35F7]=8'h00;
    mem['h35F8]=8'h00; mem['h35F9]=8'h00; mem['h35FA]=8'h00; mem['h35FB]=8'h00;
    mem['h35FC]=8'h00; mem['h35FD]=8'h00; mem['h35FE]=8'h00; mem['h35FF]=8'h00;
    mem['h3600]=8'h00; mem['h3601]=8'h00; mem['h3602]=8'h00; mem['h3603]=8'h00;
    mem['h3604]=8'h00; mem['h3605]=8'h00; mem['h3606]=8'h00; mem['h3607]=8'h00;
    mem['h3608]=8'h00; mem['h3609]=8'h00; mem['h360A]=8'h00; mem['h360B]=8'h00;
    mem['h360C]=8'h00; mem['h360D]=8'h00; mem['h360E]=8'h00; mem['h360F]=8'h00;
    mem['h3610]=8'h00; mem['h3611]=8'h00; mem['h3612]=8'h00; mem['h3613]=8'h00;
    mem['h3614]=8'h00; mem['h3615]=8'h00; mem['h3616]=8'h00; mem['h3617]=8'h00;
    mem['h3618]=8'h00; mem['h3619]=8'h00; mem['h361A]=8'h00; mem['h361B]=8'h00;
    mem['h361C]=8'h00; mem['h361D]=8'h00; mem['h361E]=8'h00; mem['h361F]=8'h00;
    mem['h3620]=8'h00; mem['h3621]=8'h00; mem['h3622]=8'h00; mem['h3623]=8'h00;
    mem['h3624]=8'h00; mem['h3625]=8'h00; mem['h3626]=8'h00; mem['h3627]=8'h00;
    mem['h3628]=8'h00; mem['h3629]=8'h00; mem['h362A]=8'h00; mem['h362B]=8'h00;
    mem['h362C]=8'h00; mem['h362D]=8'h00; mem['h362E]=8'h00; mem['h362F]=8'h00;
    mem['h3630]=8'h00; mem['h3631]=8'h00; mem['h3632]=8'h00; mem['h3633]=8'h00;
    mem['h3634]=8'h00; mem['h3635]=8'h00; mem['h3636]=8'h00; mem['h3637]=8'h00;
    mem['h3638]=8'h00; mem['h3639]=8'h00; mem['h363A]=8'h00; mem['h363B]=8'h00;
    mem['h363C]=8'h00; mem['h363D]=8'h00; mem['h363E]=8'h00; mem['h363F]=8'h00;
    mem['h3640]=8'h00; mem['h3641]=8'h00; mem['h3642]=8'h00; mem['h3643]=8'h00;
    mem['h3644]=8'h00; mem['h3645]=8'h00; mem['h3646]=8'h00; mem['h3647]=8'h00;
    mem['h3648]=8'h00; mem['h3649]=8'h00; mem['h364A]=8'h00; mem['h364B]=8'h00;
    mem['h364C]=8'h00; mem['h364D]=8'h00; mem['h364E]=8'h00; mem['h364F]=8'h00;
    mem['h3650]=8'h00; mem['h3651]=8'h00; mem['h3652]=8'h00; mem['h3653]=8'h00;
    mem['h3654]=8'h00; mem['h3655]=8'h00; mem['h3656]=8'h00; mem['h3657]=8'h00;
    mem['h3658]=8'h00; mem['h3659]=8'h00; mem['h365A]=8'h00; mem['h365B]=8'h00;
    mem['h365C]=8'h00; mem['h365D]=8'h00; mem['h365E]=8'h00; mem['h365F]=8'h00;
    mem['h3660]=8'h00; mem['h3661]=8'h00; mem['h3662]=8'h00; mem['h3663]=8'h00;
    mem['h3664]=8'h00; mem['h3665]=8'h00; mem['h3666]=8'h00; mem['h3667]=8'h00;
    mem['h3668]=8'h00; mem['h3669]=8'h00; mem['h366A]=8'h00; mem['h366B]=8'h00;
    mem['h366C]=8'h00; mem['h366D]=8'h00; mem['h366E]=8'h00; mem['h366F]=8'h00;
    mem['h3670]=8'h00; mem['h3671]=8'h00; mem['h3672]=8'h00; mem['h3673]=8'h00;
    mem['h3674]=8'h00; mem['h3675]=8'h00; mem['h3676]=8'h00; mem['h3677]=8'h00;
    mem['h3678]=8'h00; mem['h3679]=8'h00; mem['h367A]=8'h00; mem['h367B]=8'h00;
    mem['h367C]=8'h00; mem['h367D]=8'h00; mem['h367E]=8'h00; mem['h367F]=8'h00;
    mem['h3680]=8'h00; mem['h3681]=8'h00; mem['h3682]=8'h00; mem['h3683]=8'h00;
    mem['h3684]=8'h00; mem['h3685]=8'h00; mem['h3686]=8'h00; mem['h3687]=8'h00;
    mem['h3688]=8'h00; mem['h3689]=8'h00; mem['h368A]=8'h00; mem['h368B]=8'h00;
    mem['h368C]=8'h00; mem['h368D]=8'h00; mem['h368E]=8'h00; mem['h368F]=8'h00;
    mem['h3690]=8'h00; mem['h3691]=8'h00; mem['h3692]=8'h00; mem['h3693]=8'h00;
    mem['h3694]=8'h00; mem['h3695]=8'h00; mem['h3696]=8'h00; mem['h3697]=8'h00;
    mem['h3698]=8'h00; mem['h3699]=8'h00; mem['h369A]=8'h00; mem['h369B]=8'h00;
    mem['h369C]=8'h00; mem['h369D]=8'h00; mem['h369E]=8'h00; mem['h369F]=8'h00;
    mem['h36A0]=8'h00; mem['h36A1]=8'h00; mem['h36A2]=8'h00; mem['h36A3]=8'h00;
    mem['h36A4]=8'h00; mem['h36A5]=8'h00; mem['h36A6]=8'h00; mem['h36A7]=8'h00;
    mem['h36A8]=8'h00; mem['h36A9]=8'h00; mem['h36AA]=8'h00; mem['h36AB]=8'h00;
    mem['h36AC]=8'h00; mem['h36AD]=8'h00; mem['h36AE]=8'h00; mem['h36AF]=8'h00;
    mem['h36B0]=8'h00; mem['h36B1]=8'h00; mem['h36B2]=8'h00; mem['h36B3]=8'h00;
    mem['h36B4]=8'h00; mem['h36B5]=8'h00; mem['h36B6]=8'h00; mem['h36B7]=8'h00;
    mem['h36B8]=8'h00; mem['h36B9]=8'h00; mem['h36BA]=8'h00; mem['h36BB]=8'h00;
    mem['h36BC]=8'h00; mem['h36BD]=8'h00; mem['h36BE]=8'h00; mem['h36BF]=8'h00;
    mem['h36C0]=8'h00; mem['h36C1]=8'h00; mem['h36C2]=8'h00; mem['h36C3]=8'h00;
    mem['h36C4]=8'h00; mem['h36C5]=8'h00; mem['h36C6]=8'h00; mem['h36C7]=8'h00;
    mem['h36C8]=8'h00; mem['h36C9]=8'h00; mem['h36CA]=8'h00; mem['h36CB]=8'h00;
    mem['h36CC]=8'h00; mem['h36CD]=8'h00; mem['h36CE]=8'h00; mem['h36CF]=8'h00;
    mem['h36D0]=8'h00; mem['h36D1]=8'h00; mem['h36D2]=8'h00; mem['h36D3]=8'h00;
    mem['h36D4]=8'h00; mem['h36D5]=8'h00; mem['h36D6]=8'h00; mem['h36D7]=8'h00;
    mem['h36D8]=8'h00; mem['h36D9]=8'h00; mem['h36DA]=8'h00; mem['h36DB]=8'h00;
    mem['h36DC]=8'h00; mem['h36DD]=8'h00; mem['h36DE]=8'h00; mem['h36DF]=8'h00;
    mem['h36E0]=8'h00; mem['h36E1]=8'h00; mem['h36E2]=8'h00; mem['h36E3]=8'h00;
    mem['h36E4]=8'h00; mem['h36E5]=8'h00; mem['h36E6]=8'h00; mem['h36E7]=8'h00;
    mem['h36E8]=8'h00; mem['h36E9]=8'h00; mem['h36EA]=8'h00; mem['h36EB]=8'h00;
    mem['h36EC]=8'h00; mem['h36ED]=8'h00; mem['h36EE]=8'h00; mem['h36EF]=8'h00;
    mem['h36F0]=8'h00; mem['h36F1]=8'h00; mem['h36F2]=8'h00; mem['h36F3]=8'h00;
    mem['h36F4]=8'h00; mem['h36F5]=8'h00; mem['h36F6]=8'h00; mem['h36F7]=8'h00;
    mem['h36F8]=8'h00; mem['h36F9]=8'h00; mem['h36FA]=8'h00; mem['h36FB]=8'h00;
    mem['h36FC]=8'h00; mem['h36FD]=8'h00; mem['h36FE]=8'h00; mem['h36FF]=8'h00;
    mem['h3700]=8'h00; mem['h3701]=8'h00; mem['h3702]=8'h00; mem['h3703]=8'h00;
    mem['h3704]=8'h00; mem['h3705]=8'h00; mem['h3706]=8'h00; mem['h3707]=8'h00;
    mem['h3708]=8'h00; mem['h3709]=8'h00; mem['h370A]=8'h00; mem['h370B]=8'h00;
    mem['h370C]=8'h00; mem['h370D]=8'h00; mem['h370E]=8'h00; mem['h370F]=8'h00;
    mem['h3710]=8'h00; mem['h3711]=8'h00; mem['h3712]=8'h00; mem['h3713]=8'h00;
    mem['h3714]=8'h00; mem['h3715]=8'h00; mem['h3716]=8'h00; mem['h3717]=8'h00;
    mem['h3718]=8'h00; mem['h3719]=8'h00; mem['h371A]=8'h00; mem['h371B]=8'h00;
    mem['h371C]=8'h00; mem['h371D]=8'h00; mem['h371E]=8'h00; mem['h371F]=8'h00;
    mem['h3720]=8'h00; mem['h3721]=8'h00; mem['h3722]=8'h00; mem['h3723]=8'h00;
    mem['h3724]=8'h00; mem['h3725]=8'h00; mem['h3726]=8'h00; mem['h3727]=8'h00;
    mem['h3728]=8'h00; mem['h3729]=8'h00; mem['h372A]=8'h00; mem['h372B]=8'h00;
    mem['h372C]=8'h00; mem['h372D]=8'h00; mem['h372E]=8'h00; mem['h372F]=8'h00;
    mem['h3730]=8'h00; mem['h3731]=8'h00; mem['h3732]=8'h00; mem['h3733]=8'h00;
    mem['h3734]=8'h00; mem['h3735]=8'h00; mem['h3736]=8'h00; mem['h3737]=8'h00;
    mem['h3738]=8'h00; mem['h3739]=8'h00; mem['h373A]=8'h00; mem['h373B]=8'h00;
    mem['h373C]=8'h00; mem['h373D]=8'h00; mem['h373E]=8'h00; mem['h373F]=8'h00;
    mem['h3740]=8'h00; mem['h3741]=8'h00; mem['h3742]=8'h00; mem['h3743]=8'h00;
    mem['h3744]=8'h00; mem['h3745]=8'h00; mem['h3746]=8'h00; mem['h3747]=8'h00;
    mem['h3748]=8'h00; mem['h3749]=8'h00; mem['h374A]=8'h00; mem['h374B]=8'h00;
    mem['h374C]=8'h00; mem['h374D]=8'h00; mem['h374E]=8'h00; mem['h374F]=8'h00;
    mem['h3750]=8'h00; mem['h3751]=8'h00; mem['h3752]=8'h00; mem['h3753]=8'h00;
    mem['h3754]=8'h00; mem['h3755]=8'h00; mem['h3756]=8'h00; mem['h3757]=8'h00;
    mem['h3758]=8'h00; mem['h3759]=8'h00; mem['h375A]=8'h00; mem['h375B]=8'h00;
    mem['h375C]=8'h00; mem['h375D]=8'h00; mem['h375E]=8'h00; mem['h375F]=8'h00;
    mem['h3760]=8'h00; mem['h3761]=8'h00; mem['h3762]=8'h00; mem['h3763]=8'h00;
    mem['h3764]=8'h00; mem['h3765]=8'h00; mem['h3766]=8'h00; mem['h3767]=8'h00;
    mem['h3768]=8'h00; mem['h3769]=8'h00; mem['h376A]=8'h00; mem['h376B]=8'h00;
    mem['h376C]=8'h00; mem['h376D]=8'h00; mem['h376E]=8'h00; mem['h376F]=8'h00;
    mem['h3770]=8'h00; mem['h3771]=8'h00; mem['h3772]=8'h00; mem['h3773]=8'h00;
    mem['h3774]=8'h00; mem['h3775]=8'h00; mem['h3776]=8'h00; mem['h3777]=8'h00;
    mem['h3778]=8'h00; mem['h3779]=8'h00; mem['h377A]=8'h00; mem['h377B]=8'h00;
    mem['h377C]=8'h00; mem['h377D]=8'h00; mem['h377E]=8'h00; mem['h377F]=8'h00;
    mem['h3780]=8'h00; mem['h3781]=8'h00; mem['h3782]=8'h00; mem['h3783]=8'h00;
    mem['h3784]=8'h00; mem['h3785]=8'h00; mem['h3786]=8'h00; mem['h3787]=8'h00;
    mem['h3788]=8'h00; mem['h3789]=8'h00; mem['h378A]=8'h00; mem['h378B]=8'h00;
    mem['h378C]=8'h00; mem['h378D]=8'h00; mem['h378E]=8'h00; mem['h378F]=8'h00;
    mem['h3790]=8'h00; mem['h3791]=8'h00; mem['h3792]=8'h00; mem['h3793]=8'h00;
    mem['h3794]=8'h00; mem['h3795]=8'h00; mem['h3796]=8'h00; mem['h3797]=8'h00;
    mem['h3798]=8'h00; mem['h3799]=8'h00; mem['h379A]=8'h00; mem['h379B]=8'h00;
    mem['h379C]=8'h00; mem['h379D]=8'h00; mem['h379E]=8'h00; mem['h379F]=8'h00;
    mem['h37A0]=8'h00; mem['h37A1]=8'h00; mem['h37A2]=8'h00; mem['h37A3]=8'h00;
    mem['h37A4]=8'h00; mem['h37A5]=8'h00; mem['h37A6]=8'h00; mem['h37A7]=8'h00;
    mem['h37A8]=8'h00; mem['h37A9]=8'h00; mem['h37AA]=8'h00; mem['h37AB]=8'h00;
    mem['h37AC]=8'h00; mem['h37AD]=8'h00; mem['h37AE]=8'h00; mem['h37AF]=8'h00;
    mem['h37B0]=8'h00; mem['h37B1]=8'h00; mem['h37B2]=8'h00; mem['h37B3]=8'h00;
    mem['h37B4]=8'h00; mem['h37B5]=8'h00; mem['h37B6]=8'h00; mem['h37B7]=8'h00;
    mem['h37B8]=8'h00; mem['h37B9]=8'h00; mem['h37BA]=8'h00; mem['h37BB]=8'h00;
    mem['h37BC]=8'h00; mem['h37BD]=8'h00; mem['h37BE]=8'h00; mem['h37BF]=8'h00;
    mem['h37C0]=8'h00; mem['h37C1]=8'h00; mem['h37C2]=8'h00; mem['h37C3]=8'h00;
    mem['h37C4]=8'h00; mem['h37C5]=8'h00; mem['h37C6]=8'h00; mem['h37C7]=8'h00;
    mem['h37C8]=8'h00; mem['h37C9]=8'h00; mem['h37CA]=8'h00; mem['h37CB]=8'h00;
    mem['h37CC]=8'h00; mem['h37CD]=8'h00; mem['h37CE]=8'h00; mem['h37CF]=8'h00;
    mem['h37D0]=8'h00; mem['h37D1]=8'h00; mem['h37D2]=8'h00; mem['h37D3]=8'h00;
    mem['h37D4]=8'h00; mem['h37D5]=8'h00; mem['h37D6]=8'h00; mem['h37D7]=8'h00;
    mem['h37D8]=8'h00; mem['h37D9]=8'h00; mem['h37DA]=8'h00; mem['h37DB]=8'h00;
    mem['h37DC]=8'h00; mem['h37DD]=8'h00; mem['h37DE]=8'h00; mem['h37DF]=8'h00;
    mem['h37E0]=8'h00; mem['h37E1]=8'h00; mem['h37E2]=8'h00; mem['h37E3]=8'h00;
    mem['h37E4]=8'h00; mem['h37E5]=8'h00; mem['h37E6]=8'h00; mem['h37E7]=8'h00;
    mem['h37E8]=8'h00; mem['h37E9]=8'h00; mem['h37EA]=8'h00; mem['h37EB]=8'h00;
    mem['h37EC]=8'h00; mem['h37ED]=8'h00; mem['h37EE]=8'h00; mem['h37EF]=8'h00;
    mem['h37F0]=8'h00; mem['h37F1]=8'h00; mem['h37F2]=8'h00; mem['h37F3]=8'h00;
    mem['h37F4]=8'h00; mem['h37F5]=8'h00; mem['h37F6]=8'h00; mem['h37F7]=8'h00;
    mem['h37F8]=8'h00; mem['h37F9]=8'h00; mem['h37FA]=8'h00; mem['h37FB]=8'h00;
    mem['h37FC]=8'h00; mem['h37FD]=8'h00; mem['h37FE]=8'h00; mem['h37FF]=8'h00;
    mem['h3800]=8'h00; mem['h3801]=8'h00; mem['h3802]=8'h00; mem['h3803]=8'h00;
    mem['h3804]=8'h00; mem['h3805]=8'h00; mem['h3806]=8'h00; mem['h3807]=8'h00;
    mem['h3808]=8'h00; mem['h3809]=8'h00; mem['h380A]=8'h00; mem['h380B]=8'h00;
    mem['h380C]=8'h00; mem['h380D]=8'h00; mem['h380E]=8'h00; mem['h380F]=8'h00;
    mem['h3810]=8'h00; mem['h3811]=8'h00; mem['h3812]=8'h00; mem['h3813]=8'h00;
    mem['h3814]=8'h00; mem['h3815]=8'h00; mem['h3816]=8'h00; mem['h3817]=8'h00;
    mem['h3818]=8'h00; mem['h3819]=8'h00; mem['h381A]=8'h00; mem['h381B]=8'h00;
    mem['h381C]=8'h00; mem['h381D]=8'h00; mem['h381E]=8'h00; mem['h381F]=8'h00;
    mem['h3820]=8'h00; mem['h3821]=8'h00; mem['h3822]=8'h00; mem['h3823]=8'h00;
    mem['h3824]=8'h00; mem['h3825]=8'h00; mem['h3826]=8'h00; mem['h3827]=8'h00;
    mem['h3828]=8'h00; mem['h3829]=8'h00; mem['h382A]=8'h00; mem['h382B]=8'h00;
    mem['h382C]=8'h00; mem['h382D]=8'h00; mem['h382E]=8'h00; mem['h382F]=8'h00;
    mem['h3830]=8'h00; mem['h3831]=8'h00; mem['h3832]=8'h00; mem['h3833]=8'h00;
    mem['h3834]=8'h00; mem['h3835]=8'h00; mem['h3836]=8'h00; mem['h3837]=8'h00;
    mem['h3838]=8'h00; mem['h3839]=8'h00; mem['h383A]=8'h00; mem['h383B]=8'h00;
    mem['h383C]=8'h00; mem['h383D]=8'h00; mem['h383E]=8'h00; mem['h383F]=8'h00;
    mem['h3840]=8'h00; mem['h3841]=8'h00; mem['h3842]=8'h00; mem['h3843]=8'h00;
    mem['h3844]=8'h00; mem['h3845]=8'h00; mem['h3846]=8'h00; mem['h3847]=8'h00;
    mem['h3848]=8'h00; mem['h3849]=8'h00; mem['h384A]=8'h00; mem['h384B]=8'h00;
    mem['h384C]=8'h00; mem['h384D]=8'h00; mem['h384E]=8'h00; mem['h384F]=8'h00;
    mem['h3850]=8'h00; mem['h3851]=8'h00; mem['h3852]=8'h00; mem['h3853]=8'h00;
    mem['h3854]=8'h00; mem['h3855]=8'h00; mem['h3856]=8'h00; mem['h3857]=8'h00;
    mem['h3858]=8'h00; mem['h3859]=8'h00; mem['h385A]=8'h00; mem['h385B]=8'h00;
    mem['h385C]=8'h00; mem['h385D]=8'h00; mem['h385E]=8'h00; mem['h385F]=8'h00;
    mem['h3860]=8'h00; mem['h3861]=8'h00; mem['h3862]=8'h00; mem['h3863]=8'h00;
    mem['h3864]=8'h00; mem['h3865]=8'h00; mem['h3866]=8'h00; mem['h3867]=8'h00;
    mem['h3868]=8'h00; mem['h3869]=8'h00; mem['h386A]=8'h00; mem['h386B]=8'h00;
    mem['h386C]=8'h00; mem['h386D]=8'h00; mem['h386E]=8'h00; mem['h386F]=8'h00;
    mem['h3870]=8'h00; mem['h3871]=8'h00; mem['h3872]=8'h00; mem['h3873]=8'h00;
    mem['h3874]=8'h00; mem['h3875]=8'h00; mem['h3876]=8'h00; mem['h3877]=8'h00;
    mem['h3878]=8'h00; mem['h3879]=8'h00; mem['h387A]=8'h00; mem['h387B]=8'h00;
    mem['h387C]=8'h00; mem['h387D]=8'h00; mem['h387E]=8'h00; mem['h387F]=8'h00;
    mem['h3880]=8'h00; mem['h3881]=8'h00; mem['h3882]=8'h00; mem['h3883]=8'h00;
    mem['h3884]=8'h00; mem['h3885]=8'h00; mem['h3886]=8'h00; mem['h3887]=8'h00;
    mem['h3888]=8'h00; mem['h3889]=8'h00; mem['h388A]=8'h00; mem['h388B]=8'h00;
    mem['h388C]=8'h00; mem['h388D]=8'h00; mem['h388E]=8'h00; mem['h388F]=8'h00;
    mem['h3890]=8'h00; mem['h3891]=8'h00; mem['h3892]=8'h00; mem['h3893]=8'h00;
    mem['h3894]=8'h00; mem['h3895]=8'h00; mem['h3896]=8'h00; mem['h3897]=8'h00;
    mem['h3898]=8'h00; mem['h3899]=8'h00; mem['h389A]=8'h00; mem['h389B]=8'h00;
    mem['h389C]=8'h00; mem['h389D]=8'h00; mem['h389E]=8'h00; mem['h389F]=8'h00;
    mem['h38A0]=8'h00; mem['h38A1]=8'h00; mem['h38A2]=8'h00; mem['h38A3]=8'h00;
    mem['h38A4]=8'h00; mem['h38A5]=8'h00; mem['h38A6]=8'h00; mem['h38A7]=8'h00;
    mem['h38A8]=8'h00; mem['h38A9]=8'h00; mem['h38AA]=8'h00; mem['h38AB]=8'h00;
    mem['h38AC]=8'h00; mem['h38AD]=8'h00; mem['h38AE]=8'h00; mem['h38AF]=8'h00;
    mem['h38B0]=8'h00; mem['h38B1]=8'h00; mem['h38B2]=8'h00; mem['h38B3]=8'h00;
    mem['h38B4]=8'h00; mem['h38B5]=8'h00; mem['h38B6]=8'h00; mem['h38B7]=8'h00;
    mem['h38B8]=8'h00; mem['h38B9]=8'h00; mem['h38BA]=8'h00; mem['h38BB]=8'h00;
    mem['h38BC]=8'h00; mem['h38BD]=8'h00; mem['h38BE]=8'h00; mem['h38BF]=8'h00;
    mem['h38C0]=8'h00; mem['h38C1]=8'h00; mem['h38C2]=8'h00; mem['h38C3]=8'h00;
    mem['h38C4]=8'h00; mem['h38C5]=8'h00; mem['h38C6]=8'h00; mem['h38C7]=8'h00;
    mem['h38C8]=8'h00; mem['h38C9]=8'h00; mem['h38CA]=8'h00; mem['h38CB]=8'h00;
    mem['h38CC]=8'h00; mem['h38CD]=8'h00; mem['h38CE]=8'h00; mem['h38CF]=8'h00;
    mem['h38D0]=8'h00; mem['h38D1]=8'h00; mem['h38D2]=8'h00; mem['h38D3]=8'h00;
    mem['h38D4]=8'h00; mem['h38D5]=8'h00; mem['h38D6]=8'h00; mem['h38D7]=8'h00;
    mem['h38D8]=8'h00; mem['h38D9]=8'h00; mem['h38DA]=8'h00; mem['h38DB]=8'h00;
    mem['h38DC]=8'h00; mem['h38DD]=8'h00; mem['h38DE]=8'h00; mem['h38DF]=8'h00;
    mem['h38E0]=8'h00; mem['h38E1]=8'h00; mem['h38E2]=8'h00; mem['h38E3]=8'h00;
    mem['h38E4]=8'h00; mem['h38E5]=8'h00; mem['h38E6]=8'h00; mem['h38E7]=8'h00;
    mem['h38E8]=8'h00; mem['h38E9]=8'h00; mem['h38EA]=8'h00; mem['h38EB]=8'h00;
    mem['h38EC]=8'h00; mem['h38ED]=8'h00; mem['h38EE]=8'h00; mem['h38EF]=8'h00;
    mem['h38F0]=8'h00; mem['h38F1]=8'h00; mem['h38F2]=8'h00; mem['h38F3]=8'h00;
    mem['h38F4]=8'h00; mem['h38F5]=8'h00; mem['h38F6]=8'h00; mem['h38F7]=8'h00;
    mem['h38F8]=8'h00; mem['h38F9]=8'h00; mem['h38FA]=8'h00; mem['h38FB]=8'h00;
    mem['h38FC]=8'h00; mem['h38FD]=8'h00; mem['h38FE]=8'h00; mem['h38FF]=8'h00;
    mem['h3900]=8'h00; mem['h3901]=8'h00; mem['h3902]=8'h00; mem['h3903]=8'h00;
    mem['h3904]=8'h00; mem['h3905]=8'h00; mem['h3906]=8'h00; mem['h3907]=8'h00;
    mem['h3908]=8'h00; mem['h3909]=8'h00; mem['h390A]=8'h00; mem['h390B]=8'h00;
    mem['h390C]=8'h00; mem['h390D]=8'h00; mem['h390E]=8'h00; mem['h390F]=8'h00;
    mem['h3910]=8'h00; mem['h3911]=8'h00; mem['h3912]=8'h00; mem['h3913]=8'h00;
    mem['h3914]=8'h00; mem['h3915]=8'h00; mem['h3916]=8'h00; mem['h3917]=8'h00;
    mem['h3918]=8'h00; mem['h3919]=8'h00; mem['h391A]=8'h00; mem['h391B]=8'h00;
    mem['h391C]=8'h00; mem['h391D]=8'h00; mem['h391E]=8'h00; mem['h391F]=8'h00;
    mem['h3920]=8'h00; mem['h3921]=8'h00; mem['h3922]=8'h00; mem['h3923]=8'h00;
    mem['h3924]=8'h00; mem['h3925]=8'h00; mem['h3926]=8'h00; mem['h3927]=8'h00;
    mem['h3928]=8'h00; mem['h3929]=8'h00; mem['h392A]=8'h00; mem['h392B]=8'h00;
    mem['h392C]=8'h00; mem['h392D]=8'h00; mem['h392E]=8'h00; mem['h392F]=8'h00;
    mem['h3930]=8'h00; mem['h3931]=8'h00; mem['h3932]=8'h00; mem['h3933]=8'h00;
    mem['h3934]=8'h00; mem['h3935]=8'h00; mem['h3936]=8'h00; mem['h3937]=8'h00;
    mem['h3938]=8'h00; mem['h3939]=8'h00; mem['h393A]=8'h00; mem['h393B]=8'h00;
    mem['h393C]=8'h00; mem['h393D]=8'h00; mem['h393E]=8'h00; mem['h393F]=8'h00;
    mem['h3940]=8'h00; mem['h3941]=8'h00; mem['h3942]=8'h00; mem['h3943]=8'h00;
    mem['h3944]=8'h00; mem['h3945]=8'h00; mem['h3946]=8'h00; mem['h3947]=8'h00;
    mem['h3948]=8'h00; mem['h3949]=8'h00; mem['h394A]=8'h00; mem['h394B]=8'h00;
    mem['h394C]=8'h00; mem['h394D]=8'h00; mem['h394E]=8'h00; mem['h394F]=8'h00;
    mem['h3950]=8'h00; mem['h3951]=8'h00; mem['h3952]=8'h00; mem['h3953]=8'h00;
    mem['h3954]=8'h00; mem['h3955]=8'h00; mem['h3956]=8'h00; mem['h3957]=8'h00;
    mem['h3958]=8'h00; mem['h3959]=8'h00; mem['h395A]=8'h00; mem['h395B]=8'h00;
    mem['h395C]=8'h00; mem['h395D]=8'h00; mem['h395E]=8'h00; mem['h395F]=8'h00;
    mem['h3960]=8'h00; mem['h3961]=8'h00; mem['h3962]=8'h00; mem['h3963]=8'h00;
    mem['h3964]=8'h00; mem['h3965]=8'h00; mem['h3966]=8'h00; mem['h3967]=8'h00;
    mem['h3968]=8'h00; mem['h3969]=8'h00; mem['h396A]=8'h00; mem['h396B]=8'h00;
    mem['h396C]=8'h00; mem['h396D]=8'h00; mem['h396E]=8'h00; mem['h396F]=8'h00;
    mem['h3970]=8'h00; mem['h3971]=8'h00; mem['h3972]=8'h00; mem['h3973]=8'h00;
    mem['h3974]=8'h00; mem['h3975]=8'h00; mem['h3976]=8'h00; mem['h3977]=8'h00;
    mem['h3978]=8'h00; mem['h3979]=8'h00; mem['h397A]=8'h00; mem['h397B]=8'h00;
    mem['h397C]=8'h00; mem['h397D]=8'h00; mem['h397E]=8'h00; mem['h397F]=8'h00;
    mem['h3980]=8'h00; mem['h3981]=8'h00; mem['h3982]=8'h00; mem['h3983]=8'h00;
    mem['h3984]=8'h00; mem['h3985]=8'h00; mem['h3986]=8'h00; mem['h3987]=8'h00;
    mem['h3988]=8'h00; mem['h3989]=8'h00; mem['h398A]=8'h00; mem['h398B]=8'h00;
    mem['h398C]=8'h00; mem['h398D]=8'h00; mem['h398E]=8'h00; mem['h398F]=8'h00;
    mem['h3990]=8'h00; mem['h3991]=8'h00; mem['h3992]=8'h00; mem['h3993]=8'h00;
    mem['h3994]=8'h00; mem['h3995]=8'h00; mem['h3996]=8'h00; mem['h3997]=8'h00;
    mem['h3998]=8'h00; mem['h3999]=8'h00; mem['h399A]=8'h00; mem['h399B]=8'h00;
    mem['h399C]=8'h00; mem['h399D]=8'h00; mem['h399E]=8'h00; mem['h399F]=8'h00;
    mem['h39A0]=8'h00; mem['h39A1]=8'h00; mem['h39A2]=8'h00; mem['h39A3]=8'h00;
    mem['h39A4]=8'h00; mem['h39A5]=8'h00; mem['h39A6]=8'h00; mem['h39A7]=8'h00;
    mem['h39A8]=8'h00; mem['h39A9]=8'h00; mem['h39AA]=8'h00; mem['h39AB]=8'h00;
    mem['h39AC]=8'h00; mem['h39AD]=8'h00; mem['h39AE]=8'h00; mem['h39AF]=8'h00;
    mem['h39B0]=8'h00; mem['h39B1]=8'h00; mem['h39B2]=8'h00; mem['h39B3]=8'h00;
    mem['h39B4]=8'h00; mem['h39B5]=8'h00; mem['h39B6]=8'h00; mem['h39B7]=8'h00;
    mem['h39B8]=8'h00; mem['h39B9]=8'h00; mem['h39BA]=8'h00; mem['h39BB]=8'h00;
    mem['h39BC]=8'h00; mem['h39BD]=8'h00; mem['h39BE]=8'h00; mem['h39BF]=8'h00;
    mem['h39C0]=8'h00; mem['h39C1]=8'h00; mem['h39C2]=8'h00; mem['h39C3]=8'h00;
    mem['h39C4]=8'h00; mem['h39C5]=8'h00; mem['h39C6]=8'h00; mem['h39C7]=8'h00;
    mem['h39C8]=8'h00; mem['h39C9]=8'h00; mem['h39CA]=8'h00; mem['h39CB]=8'h00;
    mem['h39CC]=8'h00; mem['h39CD]=8'h00; mem['h39CE]=8'h00; mem['h39CF]=8'h00;
    mem['h39D0]=8'h00; mem['h39D1]=8'h00; mem['h39D2]=8'h00; mem['h39D3]=8'h00;
    mem['h39D4]=8'h00; mem['h39D5]=8'h00; mem['h39D6]=8'h00; mem['h39D7]=8'h00;
    mem['h39D8]=8'h00; mem['h39D9]=8'h00; mem['h39DA]=8'h00; mem['h39DB]=8'h00;
    mem['h39DC]=8'h00; mem['h39DD]=8'h00; mem['h39DE]=8'h00; mem['h39DF]=8'h00;
    mem['h39E0]=8'h00; mem['h39E1]=8'h00; mem['h39E2]=8'h00; mem['h39E3]=8'h00;
    mem['h39E4]=8'h00; mem['h39E5]=8'h00; mem['h39E6]=8'h00; mem['h39E7]=8'h00;
    mem['h39E8]=8'h00; mem['h39E9]=8'h00; mem['h39EA]=8'h00; mem['h39EB]=8'h00;
    mem['h39EC]=8'h00; mem['h39ED]=8'h00; mem['h39EE]=8'h00; mem['h39EF]=8'h00;
    mem['h39F0]=8'h00; mem['h39F1]=8'h00; mem['h39F2]=8'h00; mem['h39F3]=8'h00;
    mem['h39F4]=8'h00; mem['h39F5]=8'h00; mem['h39F6]=8'h00; mem['h39F7]=8'h00;
    mem['h39F8]=8'h00; mem['h39F9]=8'h00; mem['h39FA]=8'h00; mem['h39FB]=8'h00;
    mem['h39FC]=8'h00; mem['h39FD]=8'h00; mem['h39FE]=8'h00; mem['h39FF]=8'h00;
    mem['h3A00]=8'h00; mem['h3A01]=8'h00; mem['h3A02]=8'h00; mem['h3A03]=8'h00;
    mem['h3A04]=8'h00; mem['h3A05]=8'h00; mem['h3A06]=8'h00; mem['h3A07]=8'h00;
    mem['h3A08]=8'h00; mem['h3A09]=8'h00; mem['h3A0A]=8'h00; mem['h3A0B]=8'h00;
    mem['h3A0C]=8'h00; mem['h3A0D]=8'h00; mem['h3A0E]=8'h00; mem['h3A0F]=8'h00;
    mem['h3A10]=8'h00; mem['h3A11]=8'h00; mem['h3A12]=8'h00; mem['h3A13]=8'h00;
    mem['h3A14]=8'h00; mem['h3A15]=8'h00; mem['h3A16]=8'h00; mem['h3A17]=8'h00;
    mem['h3A18]=8'h00; mem['h3A19]=8'h00; mem['h3A1A]=8'h00; mem['h3A1B]=8'h00;
    mem['h3A1C]=8'h00; mem['h3A1D]=8'h00; mem['h3A1E]=8'h00; mem['h3A1F]=8'h00;
    mem['h3A20]=8'h00; mem['h3A21]=8'h00; mem['h3A22]=8'h00; mem['h3A23]=8'h00;
    mem['h3A24]=8'h00; mem['h3A25]=8'h00; mem['h3A26]=8'h00; mem['h3A27]=8'h00;
    mem['h3A28]=8'h00; mem['h3A29]=8'h00; mem['h3A2A]=8'h00; mem['h3A2B]=8'h00;
    mem['h3A2C]=8'h00; mem['h3A2D]=8'h00; mem['h3A2E]=8'h00; mem['h3A2F]=8'h00;
    mem['h3A30]=8'h00; mem['h3A31]=8'h00; mem['h3A32]=8'h00; mem['h3A33]=8'h00;
    mem['h3A34]=8'h00; mem['h3A35]=8'h00; mem['h3A36]=8'h00; mem['h3A37]=8'h00;
    mem['h3A38]=8'h00; mem['h3A39]=8'h00; mem['h3A3A]=8'h00; mem['h3A3B]=8'h00;
    mem['h3A3C]=8'h00; mem['h3A3D]=8'h00; mem['h3A3E]=8'h00; mem['h3A3F]=8'h00;
    mem['h3A40]=8'h00; mem['h3A41]=8'h00; mem['h3A42]=8'h00; mem['h3A43]=8'h00;
    mem['h3A44]=8'h00; mem['h3A45]=8'h00; mem['h3A46]=8'h00; mem['h3A47]=8'h00;
    mem['h3A48]=8'h00; mem['h3A49]=8'h00; mem['h3A4A]=8'h00; mem['h3A4B]=8'h00;
    mem['h3A4C]=8'h00; mem['h3A4D]=8'h00; mem['h3A4E]=8'h00; mem['h3A4F]=8'h00;
    mem['h3A50]=8'h00; mem['h3A51]=8'h00; mem['h3A52]=8'h00; mem['h3A53]=8'h00;
    mem['h3A54]=8'h00; mem['h3A55]=8'h00; mem['h3A56]=8'h00; mem['h3A57]=8'h00;
    mem['h3A58]=8'h00; mem['h3A59]=8'h00; mem['h3A5A]=8'h00; mem['h3A5B]=8'h00;
    mem['h3A5C]=8'h00; mem['h3A5D]=8'h00; mem['h3A5E]=8'h00; mem['h3A5F]=8'h00;
    mem['h3A60]=8'h00; mem['h3A61]=8'h00; mem['h3A62]=8'h00; mem['h3A63]=8'h00;
    mem['h3A64]=8'h00; mem['h3A65]=8'h00; mem['h3A66]=8'h00; mem['h3A67]=8'h00;
    mem['h3A68]=8'h00; mem['h3A69]=8'h00; mem['h3A6A]=8'h00; mem['h3A6B]=8'h00;
    mem['h3A6C]=8'h00; mem['h3A6D]=8'h00; mem['h3A6E]=8'h00; mem['h3A6F]=8'h00;
    mem['h3A70]=8'h00; mem['h3A71]=8'h00; mem['h3A72]=8'h00; mem['h3A73]=8'h00;
    mem['h3A74]=8'h00; mem['h3A75]=8'h00; mem['h3A76]=8'h00; mem['h3A77]=8'h00;
    mem['h3A78]=8'h00; mem['h3A79]=8'h00; mem['h3A7A]=8'h00; mem['h3A7B]=8'h00;
    mem['h3A7C]=8'h00; mem['h3A7D]=8'h00; mem['h3A7E]=8'h00; mem['h3A7F]=8'h00;
    mem['h3A80]=8'h00; mem['h3A81]=8'h00; mem['h3A82]=8'h00; mem['h3A83]=8'h00;
    mem['h3A84]=8'h00; mem['h3A85]=8'h00; mem['h3A86]=8'h00; mem['h3A87]=8'h00;
    mem['h3A88]=8'h00; mem['h3A89]=8'h00; mem['h3A8A]=8'h00; mem['h3A8B]=8'h00;
    mem['h3A8C]=8'h00; mem['h3A8D]=8'h00; mem['h3A8E]=8'h00; mem['h3A8F]=8'h00;
    mem['h3A90]=8'h00; mem['h3A91]=8'h00; mem['h3A92]=8'h00; mem['h3A93]=8'h00;
    mem['h3A94]=8'h00; mem['h3A95]=8'h00; mem['h3A96]=8'h00; mem['h3A97]=8'h00;
    mem['h3A98]=8'h00; mem['h3A99]=8'h00; mem['h3A9A]=8'h00; mem['h3A9B]=8'h00;
    mem['h3A9C]=8'h00; mem['h3A9D]=8'h00; mem['h3A9E]=8'h00; mem['h3A9F]=8'h00;
    mem['h3AA0]=8'h00; mem['h3AA1]=8'h00; mem['h3AA2]=8'h00; mem['h3AA3]=8'h00;
    mem['h3AA4]=8'h00; mem['h3AA5]=8'h00; mem['h3AA6]=8'h00; mem['h3AA7]=8'h00;
    mem['h3AA8]=8'h00; mem['h3AA9]=8'h00; mem['h3AAA]=8'h00; mem['h3AAB]=8'h00;
    mem['h3AAC]=8'h00; mem['h3AAD]=8'h00; mem['h3AAE]=8'h00; mem['h3AAF]=8'h00;
    mem['h3AB0]=8'h00; mem['h3AB1]=8'h00; mem['h3AB2]=8'h00; mem['h3AB3]=8'h00;
    mem['h3AB4]=8'h00; mem['h3AB5]=8'h00; mem['h3AB6]=8'h00; mem['h3AB7]=8'h00;
    mem['h3AB8]=8'h00; mem['h3AB9]=8'h00; mem['h3ABA]=8'h00; mem['h3ABB]=8'h00;
    mem['h3ABC]=8'h00; mem['h3ABD]=8'h00; mem['h3ABE]=8'h00; mem['h3ABF]=8'h00;
    mem['h3AC0]=8'h00; mem['h3AC1]=8'h00; mem['h3AC2]=8'h00; mem['h3AC3]=8'h00;
    mem['h3AC4]=8'h00; mem['h3AC5]=8'h00; mem['h3AC6]=8'h00; mem['h3AC7]=8'h00;
    mem['h3AC8]=8'h00; mem['h3AC9]=8'h00; mem['h3ACA]=8'h00; mem['h3ACB]=8'h00;
    mem['h3ACC]=8'h00; mem['h3ACD]=8'h00; mem['h3ACE]=8'h00; mem['h3ACF]=8'h00;
    mem['h3AD0]=8'h00; mem['h3AD1]=8'h00; mem['h3AD2]=8'h00; mem['h3AD3]=8'h00;
    mem['h3AD4]=8'h00; mem['h3AD5]=8'h00; mem['h3AD6]=8'h00; mem['h3AD7]=8'h00;
    mem['h3AD8]=8'h00; mem['h3AD9]=8'h00; mem['h3ADA]=8'h00; mem['h3ADB]=8'h00;
    mem['h3ADC]=8'h00; mem['h3ADD]=8'h00; mem['h3ADE]=8'h00; mem['h3ADF]=8'h00;
    mem['h3AE0]=8'h00; mem['h3AE1]=8'h00; mem['h3AE2]=8'h00; mem['h3AE3]=8'h00;
    mem['h3AE4]=8'h00; mem['h3AE5]=8'h00; mem['h3AE6]=8'h00; mem['h3AE7]=8'h00;
    mem['h3AE8]=8'h00; mem['h3AE9]=8'h00; mem['h3AEA]=8'h00; mem['h3AEB]=8'h00;
    mem['h3AEC]=8'h00; mem['h3AED]=8'h00; mem['h3AEE]=8'h00; mem['h3AEF]=8'h00;
    mem['h3AF0]=8'h00; mem['h3AF1]=8'h00; mem['h3AF2]=8'h00; mem['h3AF3]=8'h00;
    mem['h3AF4]=8'h00; mem['h3AF5]=8'h00; mem['h3AF6]=8'h00; mem['h3AF7]=8'h00;
    mem['h3AF8]=8'h00; mem['h3AF9]=8'h00; mem['h3AFA]=8'h00; mem['h3AFB]=8'h00;
    mem['h3AFC]=8'h00; mem['h3AFD]=8'h00; mem['h3AFE]=8'h00; mem['h3AFF]=8'h00;
    mem['h3B00]=8'h00; mem['h3B01]=8'h00; mem['h3B02]=8'h00; mem['h3B03]=8'h00;
    mem['h3B04]=8'h00; mem['h3B05]=8'h00; mem['h3B06]=8'h00; mem['h3B07]=8'h00;
    mem['h3B08]=8'h00; mem['h3B09]=8'h00; mem['h3B0A]=8'h00; mem['h3B0B]=8'h00;
    mem['h3B0C]=8'h00; mem['h3B0D]=8'h00; mem['h3B0E]=8'h00; mem['h3B0F]=8'h00;
    mem['h3B10]=8'h00; mem['h3B11]=8'h00; mem['h3B12]=8'h00; mem['h3B13]=8'h00;
    mem['h3B14]=8'h00; mem['h3B15]=8'h00; mem['h3B16]=8'h00; mem['h3B17]=8'h00;
    mem['h3B18]=8'h00; mem['h3B19]=8'h00; mem['h3B1A]=8'h00; mem['h3B1B]=8'h00;
    mem['h3B1C]=8'h00; mem['h3B1D]=8'h00; mem['h3B1E]=8'h00; mem['h3B1F]=8'h00;
    mem['h3B20]=8'h00; mem['h3B21]=8'h00; mem['h3B22]=8'h00; mem['h3B23]=8'h00;
    mem['h3B24]=8'h00; mem['h3B25]=8'h00; mem['h3B26]=8'h00; mem['h3B27]=8'h00;
    mem['h3B28]=8'h00; mem['h3B29]=8'h00; mem['h3B2A]=8'h00; mem['h3B2B]=8'h00;
    mem['h3B2C]=8'h00; mem['h3B2D]=8'h00; mem['h3B2E]=8'h00; mem['h3B2F]=8'h00;
    mem['h3B30]=8'h00; mem['h3B31]=8'h00; mem['h3B32]=8'h00; mem['h3B33]=8'h00;
    mem['h3B34]=8'h00; mem['h3B35]=8'h00; mem['h3B36]=8'h00; mem['h3B37]=8'h00;
    mem['h3B38]=8'h00; mem['h3B39]=8'h00; mem['h3B3A]=8'h00; mem['h3B3B]=8'h00;
    mem['h3B3C]=8'h00; mem['h3B3D]=8'h00; mem['h3B3E]=8'h00; mem['h3B3F]=8'h00;
    mem['h3B40]=8'h00; mem['h3B41]=8'h00; mem['h3B42]=8'h00; mem['h3B43]=8'h00;
    mem['h3B44]=8'h00; mem['h3B45]=8'h00; mem['h3B46]=8'h00; mem['h3B47]=8'h00;
    mem['h3B48]=8'h00; mem['h3B49]=8'h00; mem['h3B4A]=8'h00; mem['h3B4B]=8'h00;
    mem['h3B4C]=8'h00; mem['h3B4D]=8'h00; mem['h3B4E]=8'h00; mem['h3B4F]=8'h00;
    mem['h3B50]=8'h00; mem['h3B51]=8'h00; mem['h3B52]=8'h00; mem['h3B53]=8'h00;
    mem['h3B54]=8'h00; mem['h3B55]=8'h00; mem['h3B56]=8'h00; mem['h3B57]=8'h00;
    mem['h3B58]=8'h00; mem['h3B59]=8'h00; mem['h3B5A]=8'h00; mem['h3B5B]=8'h00;
    mem['h3B5C]=8'h00; mem['h3B5D]=8'h00; mem['h3B5E]=8'h00; mem['h3B5F]=8'h00;
    mem['h3B60]=8'h00; mem['h3B61]=8'h00; mem['h3B62]=8'h00; mem['h3B63]=8'h00;
    mem['h3B64]=8'h00; mem['h3B65]=8'h00; mem['h3B66]=8'h00; mem['h3B67]=8'h00;
    mem['h3B68]=8'h00; mem['h3B69]=8'h00; mem['h3B6A]=8'h00; mem['h3B6B]=8'h00;
    mem['h3B6C]=8'h00; mem['h3B6D]=8'h00; mem['h3B6E]=8'h00; mem['h3B6F]=8'h00;
    mem['h3B70]=8'h00; mem['h3B71]=8'h00; mem['h3B72]=8'h00; mem['h3B73]=8'h00;
    mem['h3B74]=8'h00; mem['h3B75]=8'h00; mem['h3B76]=8'h00; mem['h3B77]=8'h00;
    mem['h3B78]=8'h00; mem['h3B79]=8'h00; mem['h3B7A]=8'h00; mem['h3B7B]=8'h00;
    mem['h3B7C]=8'h00; mem['h3B7D]=8'h00; mem['h3B7E]=8'h00; mem['h3B7F]=8'h00;
    mem['h3B80]=8'h00; mem['h3B81]=8'h00; mem['h3B82]=8'h00; mem['h3B83]=8'h00;
    mem['h3B84]=8'h00; mem['h3B85]=8'h00; mem['h3B86]=8'h00; mem['h3B87]=8'h00;
    mem['h3B88]=8'h00; mem['h3B89]=8'h00; mem['h3B8A]=8'h00; mem['h3B8B]=8'h00;
    mem['h3B8C]=8'h00; mem['h3B8D]=8'h00; mem['h3B8E]=8'h00; mem['h3B8F]=8'h00;
    mem['h3B90]=8'h00; mem['h3B91]=8'h00; mem['h3B92]=8'h00; mem['h3B93]=8'h00;
    mem['h3B94]=8'h00; mem['h3B95]=8'h00; mem['h3B96]=8'h00; mem['h3B97]=8'h00;
    mem['h3B98]=8'h00; mem['h3B99]=8'h00; mem['h3B9A]=8'h00; mem['h3B9B]=8'h00;
    mem['h3B9C]=8'h00; mem['h3B9D]=8'h00; mem['h3B9E]=8'h00; mem['h3B9F]=8'h00;
    mem['h3BA0]=8'h00; mem['h3BA1]=8'h00; mem['h3BA2]=8'h00; mem['h3BA3]=8'h00;
    mem['h3BA4]=8'h00; mem['h3BA5]=8'h00; mem['h3BA6]=8'h00; mem['h3BA7]=8'h00;
    mem['h3BA8]=8'h00; mem['h3BA9]=8'h00; mem['h3BAA]=8'h00; mem['h3BAB]=8'h00;
    mem['h3BAC]=8'h00; mem['h3BAD]=8'h00; mem['h3BAE]=8'h00; mem['h3BAF]=8'h00;
    mem['h3BB0]=8'h00; mem['h3BB1]=8'h00; mem['h3BB2]=8'h00; mem['h3BB3]=8'h00;
    mem['h3BB4]=8'h00; mem['h3BB5]=8'h00; mem['h3BB6]=8'h00; mem['h3BB7]=8'h00;
    mem['h3BB8]=8'h00; mem['h3BB9]=8'h00; mem['h3BBA]=8'h00; mem['h3BBB]=8'h00;
    mem['h3BBC]=8'h00; mem['h3BBD]=8'h00; mem['h3BBE]=8'h00; mem['h3BBF]=8'h00;
    mem['h3BC0]=8'h00; mem['h3BC1]=8'h00; mem['h3BC2]=8'h00; mem['h3BC3]=8'h00;
    mem['h3BC4]=8'h00; mem['h3BC5]=8'h00; mem['h3BC6]=8'h00; mem['h3BC7]=8'h00;
    mem['h3BC8]=8'h00; mem['h3BC9]=8'h00; mem['h3BCA]=8'h00; mem['h3BCB]=8'h00;
    mem['h3BCC]=8'h00; mem['h3BCD]=8'h00; mem['h3BCE]=8'h00; mem['h3BCF]=8'h00;
    mem['h3BD0]=8'h00; mem['h3BD1]=8'h00; mem['h3BD2]=8'h00; mem['h3BD3]=8'h00;
    mem['h3BD4]=8'h00; mem['h3BD5]=8'h00; mem['h3BD6]=8'h00; mem['h3BD7]=8'h00;
    mem['h3BD8]=8'h00; mem['h3BD9]=8'h00; mem['h3BDA]=8'h00; mem['h3BDB]=8'h00;
    mem['h3BDC]=8'h00; mem['h3BDD]=8'h00; mem['h3BDE]=8'h00; mem['h3BDF]=8'h00;
    mem['h3BE0]=8'h00; mem['h3BE1]=8'h00; mem['h3BE2]=8'h00; mem['h3BE3]=8'h00;
    mem['h3BE4]=8'h00; mem['h3BE5]=8'h00; mem['h3BE6]=8'h00; mem['h3BE7]=8'h00;
    mem['h3BE8]=8'h00; mem['h3BE9]=8'h00; mem['h3BEA]=8'h00; mem['h3BEB]=8'h00;
    mem['h3BEC]=8'h00; mem['h3BED]=8'h00; mem['h3BEE]=8'h00; mem['h3BEF]=8'h00;
    mem['h3BF0]=8'h00; mem['h3BF1]=8'h00; mem['h3BF2]=8'h00; mem['h3BF3]=8'h00;
    mem['h3BF4]=8'h00; mem['h3BF5]=8'h00; mem['h3BF6]=8'h00; mem['h3BF7]=8'h00;
    mem['h3BF8]=8'h00; mem['h3BF9]=8'h00; mem['h3BFA]=8'h00; mem['h3BFB]=8'h00;
    mem['h3BFC]=8'h00; mem['h3BFD]=8'h00; mem['h3BFE]=8'h00; mem['h3BFF]=8'h00;
    mem['h3C00]=8'h00; mem['h3C01]=8'h00; mem['h3C02]=8'h00; mem['h3C03]=8'h00;
    mem['h3C04]=8'h00; mem['h3C05]=8'h00; mem['h3C06]=8'h00; mem['h3C07]=8'h00;
    mem['h3C08]=8'h00; mem['h3C09]=8'h00; mem['h3C0A]=8'h00; mem['h3C0B]=8'h00;
    mem['h3C0C]=8'h00; mem['h3C0D]=8'h00; mem['h3C0E]=8'h00; mem['h3C0F]=8'h00;
    mem['h3C10]=8'h00; mem['h3C11]=8'h00; mem['h3C12]=8'h00; mem['h3C13]=8'h00;
    mem['h3C14]=8'h00; mem['h3C15]=8'h00; mem['h3C16]=8'h00; mem['h3C17]=8'h00;
    mem['h3C18]=8'h00; mem['h3C19]=8'h00; mem['h3C1A]=8'h00; mem['h3C1B]=8'h00;
    mem['h3C1C]=8'h00; mem['h3C1D]=8'h00; mem['h3C1E]=8'h00; mem['h3C1F]=8'h00;
    mem['h3C20]=8'h00; mem['h3C21]=8'h00; mem['h3C22]=8'h00; mem['h3C23]=8'h00;
    mem['h3C24]=8'h00; mem['h3C25]=8'h00; mem['h3C26]=8'h00; mem['h3C27]=8'h00;
    mem['h3C28]=8'h00; mem['h3C29]=8'h00; mem['h3C2A]=8'h00; mem['h3C2B]=8'h00;
    mem['h3C2C]=8'h00; mem['h3C2D]=8'h00; mem['h3C2E]=8'h00; mem['h3C2F]=8'h00;
    mem['h3C30]=8'h00; mem['h3C31]=8'h00; mem['h3C32]=8'h00; mem['h3C33]=8'h00;
    mem['h3C34]=8'h00; mem['h3C35]=8'h00; mem['h3C36]=8'h00; mem['h3C37]=8'h00;
    mem['h3C38]=8'h00; mem['h3C39]=8'h00; mem['h3C3A]=8'h00; mem['h3C3B]=8'h00;
    mem['h3C3C]=8'h00; mem['h3C3D]=8'h00; mem['h3C3E]=8'h00; mem['h3C3F]=8'h00;
    mem['h3C40]=8'h00; mem['h3C41]=8'h00; mem['h3C42]=8'h00; mem['h3C43]=8'h00;
    mem['h3C44]=8'h00; mem['h3C45]=8'h00; mem['h3C46]=8'h00; mem['h3C47]=8'h00;
    mem['h3C48]=8'h00; mem['h3C49]=8'h00; mem['h3C4A]=8'h00; mem['h3C4B]=8'h00;
    mem['h3C4C]=8'h00; mem['h3C4D]=8'h00; mem['h3C4E]=8'h00; mem['h3C4F]=8'h00;
    mem['h3C50]=8'h00; mem['h3C51]=8'h00; mem['h3C52]=8'h00; mem['h3C53]=8'h00;
    mem['h3C54]=8'h00; mem['h3C55]=8'h00; mem['h3C56]=8'h00; mem['h3C57]=8'h00;
    mem['h3C58]=8'h00; mem['h3C59]=8'h00; mem['h3C5A]=8'h00; mem['h3C5B]=8'h00;
    mem['h3C5C]=8'h00; mem['h3C5D]=8'h00; mem['h3C5E]=8'h00; mem['h3C5F]=8'h00;
    mem['h3C60]=8'h00; mem['h3C61]=8'h00; mem['h3C62]=8'h00; mem['h3C63]=8'h00;
    mem['h3C64]=8'h00; mem['h3C65]=8'h00; mem['h3C66]=8'h00; mem['h3C67]=8'h00;
    mem['h3C68]=8'h00; mem['h3C69]=8'h00; mem['h3C6A]=8'h00; mem['h3C6B]=8'h00;
    mem['h3C6C]=8'h00; mem['h3C6D]=8'h00; mem['h3C6E]=8'h00; mem['h3C6F]=8'h00;
    mem['h3C70]=8'h00; mem['h3C71]=8'h00; mem['h3C72]=8'h00; mem['h3C73]=8'h00;
    mem['h3C74]=8'h00; mem['h3C75]=8'h00; mem['h3C76]=8'h00; mem['h3C77]=8'h00;
    mem['h3C78]=8'h00; mem['h3C79]=8'h00; mem['h3C7A]=8'h00; mem['h3C7B]=8'h00;
    mem['h3C7C]=8'h00; mem['h3C7D]=8'h00; mem['h3C7E]=8'h00; mem['h3C7F]=8'h00;
    mem['h3C80]=8'h00; mem['h3C81]=8'h00; mem['h3C82]=8'h00; mem['h3C83]=8'h00;
    mem['h3C84]=8'h00; mem['h3C85]=8'h00; mem['h3C86]=8'h00; mem['h3C87]=8'h00;
    mem['h3C88]=8'h00; mem['h3C89]=8'h00; mem['h3C8A]=8'h00; mem['h3C8B]=8'h00;
    mem['h3C8C]=8'h00; mem['h3C8D]=8'h00; mem['h3C8E]=8'h00; mem['h3C8F]=8'h00;
    mem['h3C90]=8'h00; mem['h3C91]=8'h00; mem['h3C92]=8'h00; mem['h3C93]=8'h00;
    mem['h3C94]=8'h00; mem['h3C95]=8'h00; mem['h3C96]=8'h00; mem['h3C97]=8'h00;
    mem['h3C98]=8'h00; mem['h3C99]=8'h00; mem['h3C9A]=8'h00; mem['h3C9B]=8'h00;
    mem['h3C9C]=8'h00; mem['h3C9D]=8'h00; mem['h3C9E]=8'h00; mem['h3C9F]=8'h00;
    mem['h3CA0]=8'h00; mem['h3CA1]=8'h00; mem['h3CA2]=8'h00; mem['h3CA3]=8'h00;
    mem['h3CA4]=8'h00; mem['h3CA5]=8'h00; mem['h3CA6]=8'h00; mem['h3CA7]=8'h00;
    mem['h3CA8]=8'h00; mem['h3CA9]=8'h00; mem['h3CAA]=8'h00; mem['h3CAB]=8'h00;
    mem['h3CAC]=8'h00; mem['h3CAD]=8'h00; mem['h3CAE]=8'h00; mem['h3CAF]=8'h00;
    mem['h3CB0]=8'h00; mem['h3CB1]=8'h00; mem['h3CB2]=8'h00; mem['h3CB3]=8'h00;
    mem['h3CB4]=8'h00; mem['h3CB5]=8'h00; mem['h3CB6]=8'h00; mem['h3CB7]=8'h00;
    mem['h3CB8]=8'h00; mem['h3CB9]=8'h00; mem['h3CBA]=8'h00; mem['h3CBB]=8'h00;
    mem['h3CBC]=8'h00; mem['h3CBD]=8'h00; mem['h3CBE]=8'h00; mem['h3CBF]=8'h00;
    mem['h3CC0]=8'h00; mem['h3CC1]=8'h00; mem['h3CC2]=8'h00; mem['h3CC3]=8'h00;
    mem['h3CC4]=8'h00; mem['h3CC5]=8'h00; mem['h3CC6]=8'h00; mem['h3CC7]=8'h00;
    mem['h3CC8]=8'h00; mem['h3CC9]=8'h00; mem['h3CCA]=8'h00; mem['h3CCB]=8'h00;
    mem['h3CCC]=8'h00; mem['h3CCD]=8'h00; mem['h3CCE]=8'h00; mem['h3CCF]=8'h00;
    mem['h3CD0]=8'h00; mem['h3CD1]=8'h00; mem['h3CD2]=8'h00; mem['h3CD3]=8'h00;
    mem['h3CD4]=8'h00; mem['h3CD5]=8'h00; mem['h3CD6]=8'h00; mem['h3CD7]=8'h00;
    mem['h3CD8]=8'h00; mem['h3CD9]=8'h00; mem['h3CDA]=8'h00; mem['h3CDB]=8'h00;
    mem['h3CDC]=8'h00; mem['h3CDD]=8'h00; mem['h3CDE]=8'h00; mem['h3CDF]=8'h00;
    mem['h3CE0]=8'h00; mem['h3CE1]=8'h00; mem['h3CE2]=8'h00; mem['h3CE3]=8'h00;
    mem['h3CE4]=8'h00; mem['h3CE5]=8'h00; mem['h3CE6]=8'h00; mem['h3CE7]=8'h00;
    mem['h3CE8]=8'h00; mem['h3CE9]=8'h00; mem['h3CEA]=8'h00; mem['h3CEB]=8'h00;
    mem['h3CEC]=8'h00; mem['h3CED]=8'h00; mem['h3CEE]=8'h00; mem['h3CEF]=8'h00;
    mem['h3CF0]=8'h00; mem['h3CF1]=8'h00; mem['h3CF2]=8'h00; mem['h3CF3]=8'h00;
    mem['h3CF4]=8'h00; mem['h3CF5]=8'h00; mem['h3CF6]=8'h00; mem['h3CF7]=8'h00;
    mem['h3CF8]=8'h00; mem['h3CF9]=8'h00; mem['h3CFA]=8'h00; mem['h3CFB]=8'h00;
    mem['h3CFC]=8'h00; mem['h3CFD]=8'h00; mem['h3CFE]=8'h00; mem['h3CFF]=8'h00;
    mem['h3D00]=8'h00; mem['h3D01]=8'h00; mem['h3D02]=8'h00; mem['h3D03]=8'h00;
    mem['h3D04]=8'h00; mem['h3D05]=8'h00; mem['h3D06]=8'h00; mem['h3D07]=8'h00;
    mem['h3D08]=8'h00; mem['h3D09]=8'h00; mem['h3D0A]=8'h00; mem['h3D0B]=8'h00;
    mem['h3D0C]=8'h00; mem['h3D0D]=8'h00; mem['h3D0E]=8'h00; mem['h3D0F]=8'h00;
    mem['h3D10]=8'h00; mem['h3D11]=8'h00; mem['h3D12]=8'h00; mem['h3D13]=8'h00;
    mem['h3D14]=8'h00; mem['h3D15]=8'h00; mem['h3D16]=8'h00; mem['h3D17]=8'h00;
    mem['h3D18]=8'h00; mem['h3D19]=8'h00; mem['h3D1A]=8'h00; mem['h3D1B]=8'h00;
    mem['h3D1C]=8'h00; mem['h3D1D]=8'h00; mem['h3D1E]=8'h00; mem['h3D1F]=8'h00;
    mem['h3D20]=8'h00; mem['h3D21]=8'h00; mem['h3D22]=8'h00; mem['h3D23]=8'h00;
    mem['h3D24]=8'h00; mem['h3D25]=8'h00; mem['h3D26]=8'h00; mem['h3D27]=8'h00;
    mem['h3D28]=8'h00; mem['h3D29]=8'h00; mem['h3D2A]=8'h00; mem['h3D2B]=8'h00;
    mem['h3D2C]=8'h00; mem['h3D2D]=8'h00; mem['h3D2E]=8'h00; mem['h3D2F]=8'h00;
    mem['h3D30]=8'h00; mem['h3D31]=8'h00; mem['h3D32]=8'h00; mem['h3D33]=8'h00;
    mem['h3D34]=8'h00; mem['h3D35]=8'h00; mem['h3D36]=8'h00; mem['h3D37]=8'h00;
    mem['h3D38]=8'h00; mem['h3D39]=8'h00; mem['h3D3A]=8'h00; mem['h3D3B]=8'h00;
    mem['h3D3C]=8'h00; mem['h3D3D]=8'h00; mem['h3D3E]=8'h00; mem['h3D3F]=8'h00;
    mem['h3D40]=8'h00; mem['h3D41]=8'h00; mem['h3D42]=8'h00; mem['h3D43]=8'h00;
    mem['h3D44]=8'h00; mem['h3D45]=8'h00; mem['h3D46]=8'h00; mem['h3D47]=8'h00;
    mem['h3D48]=8'h00; mem['h3D49]=8'h00; mem['h3D4A]=8'h00; mem['h3D4B]=8'h00;
    mem['h3D4C]=8'h00; mem['h3D4D]=8'h00; mem['h3D4E]=8'h00; mem['h3D4F]=8'h00;
    mem['h3D50]=8'h00; mem['h3D51]=8'h00; mem['h3D52]=8'h00; mem['h3D53]=8'h00;
    mem['h3D54]=8'h00; mem['h3D55]=8'h00; mem['h3D56]=8'h00; mem['h3D57]=8'h00;
    mem['h3D58]=8'h00; mem['h3D59]=8'h00; mem['h3D5A]=8'h00; mem['h3D5B]=8'h00;
    mem['h3D5C]=8'h00; mem['h3D5D]=8'h00; mem['h3D5E]=8'h00; mem['h3D5F]=8'h00;
    mem['h3D60]=8'h00; mem['h3D61]=8'h00; mem['h3D62]=8'h00; mem['h3D63]=8'h00;
    mem['h3D64]=8'h00; mem['h3D65]=8'h00; mem['h3D66]=8'h00; mem['h3D67]=8'h00;
    mem['h3D68]=8'h00; mem['h3D69]=8'h00; mem['h3D6A]=8'h00; mem['h3D6B]=8'h00;
    mem['h3D6C]=8'h00; mem['h3D6D]=8'h00; mem['h3D6E]=8'h00; mem['h3D6F]=8'h00;
    mem['h3D70]=8'h00; mem['h3D71]=8'h00; mem['h3D72]=8'h00; mem['h3D73]=8'h00;
    mem['h3D74]=8'h00; mem['h3D75]=8'h00; mem['h3D76]=8'h00; mem['h3D77]=8'h00;
    mem['h3D78]=8'h00; mem['h3D79]=8'h00; mem['h3D7A]=8'h00; mem['h3D7B]=8'h00;
    mem['h3D7C]=8'h00; mem['h3D7D]=8'h00; mem['h3D7E]=8'h00; mem['h3D7F]=8'h00;
    mem['h3D80]=8'h00; mem['h3D81]=8'h00; mem['h3D82]=8'h00; mem['h3D83]=8'h00;
    mem['h3D84]=8'h00; mem['h3D85]=8'h00; mem['h3D86]=8'h00; mem['h3D87]=8'h00;
    mem['h3D88]=8'h00; mem['h3D89]=8'h00; mem['h3D8A]=8'h00; mem['h3D8B]=8'h00;
    mem['h3D8C]=8'h00; mem['h3D8D]=8'h00; mem['h3D8E]=8'h00; mem['h3D8F]=8'h00;
    mem['h3D90]=8'h00; mem['h3D91]=8'h00; mem['h3D92]=8'h00; mem['h3D93]=8'h00;
    mem['h3D94]=8'h00; mem['h3D95]=8'h00; mem['h3D96]=8'h00; mem['h3D97]=8'h00;
    mem['h3D98]=8'h00; mem['h3D99]=8'h00; mem['h3D9A]=8'h00; mem['h3D9B]=8'h00;
    mem['h3D9C]=8'h00; mem['h3D9D]=8'h00; mem['h3D9E]=8'h00; mem['h3D9F]=8'h00;
    mem['h3DA0]=8'h00; mem['h3DA1]=8'h00; mem['h3DA2]=8'h00; mem['h3DA3]=8'h00;
    mem['h3DA4]=8'h00; mem['h3DA5]=8'h00; mem['h3DA6]=8'h00; mem['h3DA7]=8'h00;
    mem['h3DA8]=8'h00; mem['h3DA9]=8'h00; mem['h3DAA]=8'h00; mem['h3DAB]=8'h00;
    mem['h3DAC]=8'h00; mem['h3DAD]=8'h00; mem['h3DAE]=8'h00; mem['h3DAF]=8'h00;
    mem['h3DB0]=8'h00; mem['h3DB1]=8'h00; mem['h3DB2]=8'h00; mem['h3DB3]=8'h00;
    mem['h3DB4]=8'h00; mem['h3DB5]=8'h00; mem['h3DB6]=8'h00; mem['h3DB7]=8'h00;
    mem['h3DB8]=8'h00; mem['h3DB9]=8'h00; mem['h3DBA]=8'h00; mem['h3DBB]=8'h00;
    mem['h3DBC]=8'h00; mem['h3DBD]=8'h00; mem['h3DBE]=8'h00; mem['h3DBF]=8'h00;
    mem['h3DC0]=8'h00; mem['h3DC1]=8'h00; mem['h3DC2]=8'h00; mem['h3DC3]=8'h00;
    mem['h3DC4]=8'h00; mem['h3DC5]=8'h00; mem['h3DC6]=8'h00; mem['h3DC7]=8'h00;
    mem['h3DC8]=8'h00; mem['h3DC9]=8'h00; mem['h3DCA]=8'h00; mem['h3DCB]=8'h00;
    mem['h3DCC]=8'h00; mem['h3DCD]=8'h00; mem['h3DCE]=8'h00; mem['h3DCF]=8'h00;
    mem['h3DD0]=8'h00; mem['h3DD1]=8'h00; mem['h3DD2]=8'h00; mem['h3DD3]=8'h00;
    mem['h3DD4]=8'h00; mem['h3DD5]=8'h00; mem['h3DD6]=8'h00; mem['h3DD7]=8'h00;
    mem['h3DD8]=8'h00; mem['h3DD9]=8'h00; mem['h3DDA]=8'h00; mem['h3DDB]=8'h00;
    mem['h3DDC]=8'h00; mem['h3DDD]=8'h00; mem['h3DDE]=8'h00; mem['h3DDF]=8'h00;
    mem['h3DE0]=8'h00; mem['h3DE1]=8'h00; mem['h3DE2]=8'h00; mem['h3DE3]=8'h00;
    mem['h3DE4]=8'h00; mem['h3DE5]=8'h00; mem['h3DE6]=8'h00; mem['h3DE7]=8'h00;
    mem['h3DE8]=8'h00; mem['h3DE9]=8'h00; mem['h3DEA]=8'h00; mem['h3DEB]=8'h00;
    mem['h3DEC]=8'h00; mem['h3DED]=8'h00; mem['h3DEE]=8'h00; mem['h3DEF]=8'h00;
    mem['h3DF0]=8'h00; mem['h3DF1]=8'h00; mem['h3DF2]=8'h00; mem['h3DF3]=8'h00;
    mem['h3DF4]=8'h00; mem['h3DF5]=8'h00; mem['h3DF6]=8'h00; mem['h3DF7]=8'h00;
    mem['h3DF8]=8'h00; mem['h3DF9]=8'h00; mem['h3DFA]=8'h00; mem['h3DFB]=8'h00;
    mem['h3DFC]=8'h00; mem['h3DFD]=8'h00; mem['h3DFE]=8'h00; mem['h3DFF]=8'h00;
    mem['h3E00]=8'h00; mem['h3E01]=8'h00; mem['h3E02]=8'h00; mem['h3E03]=8'h00;
    mem['h3E04]=8'h00; mem['h3E05]=8'h00; mem['h3E06]=8'h00; mem['h3E07]=8'h00;
    mem['h3E08]=8'h00; mem['h3E09]=8'h00; mem['h3E0A]=8'h00; mem['h3E0B]=8'h00;
    mem['h3E0C]=8'h00; mem['h3E0D]=8'h00; mem['h3E0E]=8'h00; mem['h3E0F]=8'h00;
    mem['h3E10]=8'h00; mem['h3E11]=8'h00; mem['h3E12]=8'h00; mem['h3E13]=8'h00;
    mem['h3E14]=8'h00; mem['h3E15]=8'h00; mem['h3E16]=8'h00; mem['h3E17]=8'h00;
    mem['h3E18]=8'h00; mem['h3E19]=8'h00; mem['h3E1A]=8'h00; mem['h3E1B]=8'h00;
    mem['h3E1C]=8'h00; mem['h3E1D]=8'h00; mem['h3E1E]=8'h00; mem['h3E1F]=8'h00;
    mem['h3E20]=8'h00; mem['h3E21]=8'h00; mem['h3E22]=8'h00; mem['h3E23]=8'h00;
    mem['h3E24]=8'h00; mem['h3E25]=8'h00; mem['h3E26]=8'h00; mem['h3E27]=8'h00;
    mem['h3E28]=8'h00; mem['h3E29]=8'h00; mem['h3E2A]=8'h00; mem['h3E2B]=8'h00;
    mem['h3E2C]=8'h00; mem['h3E2D]=8'h00; mem['h3E2E]=8'h00; mem['h3E2F]=8'h00;
    mem['h3E30]=8'h00; mem['h3E31]=8'h00; mem['h3E32]=8'h00; mem['h3E33]=8'h00;
    mem['h3E34]=8'h00; mem['h3E35]=8'h00; mem['h3E36]=8'h00; mem['h3E37]=8'h00;
    mem['h3E38]=8'h00; mem['h3E39]=8'h00; mem['h3E3A]=8'h00; mem['h3E3B]=8'h00;
    mem['h3E3C]=8'h00; mem['h3E3D]=8'h00; mem['h3E3E]=8'h00; mem['h3E3F]=8'h00;
    mem['h3E40]=8'h00; mem['h3E41]=8'h00; mem['h3E42]=8'h00; mem['h3E43]=8'h00;
    mem['h3E44]=8'h00; mem['h3E45]=8'h00; mem['h3E46]=8'h00; mem['h3E47]=8'h00;
    mem['h3E48]=8'h00; mem['h3E49]=8'h00; mem['h3E4A]=8'h00; mem['h3E4B]=8'h00;
    mem['h3E4C]=8'h00; mem['h3E4D]=8'h00; mem['h3E4E]=8'h00; mem['h3E4F]=8'h00;
    mem['h3E50]=8'h00; mem['h3E51]=8'h00; mem['h3E52]=8'h00; mem['h3E53]=8'h00;
    mem['h3E54]=8'h00; mem['h3E55]=8'h00; mem['h3E56]=8'h00; mem['h3E57]=8'h00;
    mem['h3E58]=8'h00; mem['h3E59]=8'h00; mem['h3E5A]=8'h00; mem['h3E5B]=8'h00;
    mem['h3E5C]=8'h00; mem['h3E5D]=8'h00; mem['h3E5E]=8'h00; mem['h3E5F]=8'h00;
    mem['h3E60]=8'h00; mem['h3E61]=8'h00; mem['h3E62]=8'h00; mem['h3E63]=8'h00;
    mem['h3E64]=8'h00; mem['h3E65]=8'h00; mem['h3E66]=8'h00; mem['h3E67]=8'h00;
    mem['h3E68]=8'h00; mem['h3E69]=8'h00; mem['h3E6A]=8'h00; mem['h3E6B]=8'h00;
    mem['h3E6C]=8'h00; mem['h3E6D]=8'h00; mem['h3E6E]=8'h00; mem['h3E6F]=8'h00;
    mem['h3E70]=8'h00; mem['h3E71]=8'h00; mem['h3E72]=8'h00; mem['h3E73]=8'h00;
    mem['h3E74]=8'h00; mem['h3E75]=8'h00; mem['h3E76]=8'h00; mem['h3E77]=8'h00;
    mem['h3E78]=8'h00; mem['h3E79]=8'h00; mem['h3E7A]=8'h00; mem['h3E7B]=8'h00;
    mem['h3E7C]=8'h00; mem['h3E7D]=8'h00; mem['h3E7E]=8'h00; mem['h3E7F]=8'h00;
    mem['h3E80]=8'h00; mem['h3E81]=8'h00; mem['h3E82]=8'h00; mem['h3E83]=8'h00;
    mem['h3E84]=8'h00; mem['h3E85]=8'h00; mem['h3E86]=8'h00; mem['h3E87]=8'h00;
    mem['h3E88]=8'h00; mem['h3E89]=8'h00; mem['h3E8A]=8'h00; mem['h3E8B]=8'h00;
    mem['h3E8C]=8'h00; mem['h3E8D]=8'h00; mem['h3E8E]=8'h00; mem['h3E8F]=8'h00;
    mem['h3E90]=8'h00; mem['h3E91]=8'h00; mem['h3E92]=8'h00; mem['h3E93]=8'h00;
    mem['h3E94]=8'h00; mem['h3E95]=8'h00; mem['h3E96]=8'h00; mem['h3E97]=8'h00;
    mem['h3E98]=8'h00; mem['h3E99]=8'h00; mem['h3E9A]=8'h00; mem['h3E9B]=8'h00;
    mem['h3E9C]=8'h00; mem['h3E9D]=8'h00; mem['h3E9E]=8'h00; mem['h3E9F]=8'h00;
    mem['h3EA0]=8'h00; mem['h3EA1]=8'h00; mem['h3EA2]=8'h00; mem['h3EA3]=8'h00;
    mem['h3EA4]=8'h00; mem['h3EA5]=8'h00; mem['h3EA6]=8'h00; mem['h3EA7]=8'h00;
    mem['h3EA8]=8'h00; mem['h3EA9]=8'h00; mem['h3EAA]=8'h00; mem['h3EAB]=8'h00;
    mem['h3EAC]=8'h00; mem['h3EAD]=8'h00; mem['h3EAE]=8'h00; mem['h3EAF]=8'h00;
    mem['h3EB0]=8'h00; mem['h3EB1]=8'h00; mem['h3EB2]=8'h00; mem['h3EB3]=8'h00;
    mem['h3EB4]=8'h00; mem['h3EB5]=8'h00; mem['h3EB6]=8'h00; mem['h3EB7]=8'h00;
    mem['h3EB8]=8'h00; mem['h3EB9]=8'h00; mem['h3EBA]=8'h00; mem['h3EBB]=8'h00;
    mem['h3EBC]=8'h00; mem['h3EBD]=8'h00; mem['h3EBE]=8'h00; mem['h3EBF]=8'h00;
    mem['h3EC0]=8'h00; mem['h3EC1]=8'h00; mem['h3EC2]=8'h00; mem['h3EC3]=8'h00;
    mem['h3EC4]=8'h00; mem['h3EC5]=8'h00; mem['h3EC6]=8'h00; mem['h3EC7]=8'h00;
    mem['h3EC8]=8'h00; mem['h3EC9]=8'h00; mem['h3ECA]=8'h00; mem['h3ECB]=8'h00;
    mem['h3ECC]=8'h00; mem['h3ECD]=8'h00; mem['h3ECE]=8'h00; mem['h3ECF]=8'h00;
    mem['h3ED0]=8'h00; mem['h3ED1]=8'h00; mem['h3ED2]=8'h00; mem['h3ED3]=8'h00;
    mem['h3ED4]=8'h00; mem['h3ED5]=8'h00; mem['h3ED6]=8'h00; mem['h3ED7]=8'h00;
    mem['h3ED8]=8'h00; mem['h3ED9]=8'h00; mem['h3EDA]=8'h00; mem['h3EDB]=8'h00;
    mem['h3EDC]=8'h00; mem['h3EDD]=8'h00; mem['h3EDE]=8'h00; mem['h3EDF]=8'h00;
    mem['h3EE0]=8'h00; mem['h3EE1]=8'h00; mem['h3EE2]=8'h00; mem['h3EE3]=8'h00;
    mem['h3EE4]=8'h00; mem['h3EE5]=8'h00; mem['h3EE6]=8'h00; mem['h3EE7]=8'h00;
    mem['h3EE8]=8'h00; mem['h3EE9]=8'h00; mem['h3EEA]=8'h00; mem['h3EEB]=8'h00;
    mem['h3EEC]=8'h00; mem['h3EED]=8'h00; mem['h3EEE]=8'h00; mem['h3EEF]=8'h00;
    mem['h3EF0]=8'h00; mem['h3EF1]=8'h00; mem['h3EF2]=8'h00; mem['h3EF3]=8'h00;
    mem['h3EF4]=8'h00; mem['h3EF5]=8'h00; mem['h3EF6]=8'h00; mem['h3EF7]=8'h00;
    mem['h3EF8]=8'h00; mem['h3EF9]=8'h00; mem['h3EFA]=8'h00; mem['h3EFB]=8'h00;
    mem['h3EFC]=8'h00; mem['h3EFD]=8'h00; mem['h3EFE]=8'h00; mem['h3EFF]=8'h00;
    mem['h3F00]=8'h00; mem['h3F01]=8'h00; mem['h3F02]=8'h00; mem['h3F03]=8'h00;
    mem['h3F04]=8'h00; mem['h3F05]=8'h00; mem['h3F06]=8'h00; mem['h3F07]=8'h00;
    mem['h3F08]=8'h00; mem['h3F09]=8'h00; mem['h3F0A]=8'h00; mem['h3F0B]=8'h00;
    mem['h3F0C]=8'h00; mem['h3F0D]=8'h00; mem['h3F0E]=8'h00; mem['h3F0F]=8'h00;
    mem['h3F10]=8'h00; mem['h3F11]=8'h00; mem['h3F12]=8'h00; mem['h3F13]=8'h00;
    mem['h3F14]=8'h00; mem['h3F15]=8'h00; mem['h3F16]=8'h00; mem['h3F17]=8'h00;
    mem['h3F18]=8'h00; mem['h3F19]=8'h00; mem['h3F1A]=8'h00; mem['h3F1B]=8'h00;
    mem['h3F1C]=8'h00; mem['h3F1D]=8'h00; mem['h3F1E]=8'h00; mem['h3F1F]=8'h00;
    mem['h3F20]=8'h00; mem['h3F21]=8'h00; mem['h3F22]=8'h00; mem['h3F23]=8'h00;
    mem['h3F24]=8'h00; mem['h3F25]=8'h00; mem['h3F26]=8'h00; mem['h3F27]=8'h00;
    mem['h3F28]=8'h00; mem['h3F29]=8'h00; mem['h3F2A]=8'h00; mem['h3F2B]=8'h00;
    mem['h3F2C]=8'h00; mem['h3F2D]=8'h00; mem['h3F2E]=8'h00; mem['h3F2F]=8'h00;
    mem['h3F30]=8'h00; mem['h3F31]=8'h00; mem['h3F32]=8'h00; mem['h3F33]=8'h00;
    mem['h3F34]=8'h00; mem['h3F35]=8'h00; mem['h3F36]=8'h00; mem['h3F37]=8'h00;
    mem['h3F38]=8'h00; mem['h3F39]=8'h00; mem['h3F3A]=8'h00; mem['h3F3B]=8'h00;
    mem['h3F3C]=8'h00; mem['h3F3D]=8'h00; mem['h3F3E]=8'h00; mem['h3F3F]=8'h00;
    mem['h3F40]=8'h00; mem['h3F41]=8'h00; mem['h3F42]=8'h00; mem['h3F43]=8'h00;
    mem['h3F44]=8'h00; mem['h3F45]=8'h00; mem['h3F46]=8'h00; mem['h3F47]=8'h00;
    mem['h3F48]=8'h00; mem['h3F49]=8'h00; mem['h3F4A]=8'h00; mem['h3F4B]=8'h00;
    mem['h3F4C]=8'h00; mem['h3F4D]=8'h00; mem['h3F4E]=8'h00; mem['h3F4F]=8'h00;
    mem['h3F50]=8'h00; mem['h3F51]=8'h00; mem['h3F52]=8'h00; mem['h3F53]=8'h00;
    mem['h3F54]=8'h00; mem['h3F55]=8'h00; mem['h3F56]=8'h00; mem['h3F57]=8'h00;
    mem['h3F58]=8'h00; mem['h3F59]=8'h00; mem['h3F5A]=8'h00; mem['h3F5B]=8'h00;
    mem['h3F5C]=8'h00; mem['h3F5D]=8'h00; mem['h3F5E]=8'h00; mem['h3F5F]=8'h00;
    mem['h3F60]=8'h00; mem['h3F61]=8'h00; mem['h3F62]=8'h00; mem['h3F63]=8'h00;
    mem['h3F64]=8'h00; mem['h3F65]=8'h00; mem['h3F66]=8'h00; mem['h3F67]=8'h00;
    mem['h3F68]=8'h00; mem['h3F69]=8'h00; mem['h3F6A]=8'h00; mem['h3F6B]=8'h00;
    mem['h3F6C]=8'h00; mem['h3F6D]=8'h00; mem['h3F6E]=8'h00; mem['h3F6F]=8'h00;
    mem['h3F70]=8'h00; mem['h3F71]=8'h00; mem['h3F72]=8'h00; mem['h3F73]=8'h00;
    mem['h3F74]=8'h00; mem['h3F75]=8'h00; mem['h3F76]=8'h00; mem['h3F77]=8'h00;
    mem['h3F78]=8'h00; mem['h3F79]=8'h00; mem['h3F7A]=8'h00; mem['h3F7B]=8'h00;
    mem['h3F7C]=8'h00; mem['h3F7D]=8'h00; mem['h3F7E]=8'h00; mem['h3F7F]=8'h00;
    mem['h3F80]=8'h00; mem['h3F81]=8'h00; mem['h3F82]=8'h00; mem['h3F83]=8'h00;
    mem['h3F84]=8'h00; mem['h3F85]=8'h00; mem['h3F86]=8'h00; mem['h3F87]=8'h00;
    mem['h3F88]=8'h00; mem['h3F89]=8'h00; mem['h3F8A]=8'h00; mem['h3F8B]=8'h00;
    mem['h3F8C]=8'h00; mem['h3F8D]=8'h00; mem['h3F8E]=8'h00; mem['h3F8F]=8'h00;
    mem['h3F90]=8'h00; mem['h3F91]=8'h00; mem['h3F92]=8'h00; mem['h3F93]=8'h00;
    mem['h3F94]=8'h00; mem['h3F95]=8'h00; mem['h3F96]=8'h00; mem['h3F97]=8'h00;
    mem['h3F98]=8'h00; mem['h3F99]=8'h00; mem['h3F9A]=8'h00; mem['h3F9B]=8'h00;
    mem['h3F9C]=8'h00; mem['h3F9D]=8'h00; mem['h3F9E]=8'h00; mem['h3F9F]=8'h00;
    mem['h3FA0]=8'h00; mem['h3FA1]=8'h00; mem['h3FA2]=8'h00; mem['h3FA3]=8'h00;
    mem['h3FA4]=8'h00; mem['h3FA5]=8'h00; mem['h3FA6]=8'h00; mem['h3FA7]=8'h00;
    mem['h3FA8]=8'h00; mem['h3FA9]=8'h00; mem['h3FAA]=8'h00; mem['h3FAB]=8'h00;
    mem['h3FAC]=8'h00; mem['h3FAD]=8'h00; mem['h3FAE]=8'h00; mem['h3FAF]=8'h00;
    mem['h3FB0]=8'h00; mem['h3FB1]=8'h00; mem['h3FB2]=8'h00; mem['h3FB3]=8'h00;
    mem['h3FB4]=8'h00; mem['h3FB5]=8'h00; mem['h3FB6]=8'h00; mem['h3FB7]=8'h00;
    mem['h3FB8]=8'h00; mem['h3FB9]=8'h00; mem['h3FBA]=8'h00; mem['h3FBB]=8'h00;
    mem['h3FBC]=8'h00; mem['h3FBD]=8'h00; mem['h3FBE]=8'h00; mem['h3FBF]=8'h00;
    mem['h3FC0]=8'h00; mem['h3FC1]=8'h00; mem['h3FC2]=8'h00; mem['h3FC3]=8'h00;
    mem['h3FC4]=8'h00; mem['h3FC5]=8'h00; mem['h3FC6]=8'h00; mem['h3FC7]=8'h00;
    mem['h3FC8]=8'h00; mem['h3FC9]=8'h00; mem['h3FCA]=8'h00; mem['h3FCB]=8'h00;
    mem['h3FCC]=8'h00; mem['h3FCD]=8'h00; mem['h3FCE]=8'h00; mem['h3FCF]=8'h00;
    mem['h3FD0]=8'h00; mem['h3FD1]=8'h00; mem['h3FD2]=8'h00; mem['h3FD3]=8'h00;
    mem['h3FD4]=8'h00; mem['h3FD5]=8'h00; mem['h3FD6]=8'h00; mem['h3FD7]=8'h00;
    mem['h3FD8]=8'h00; mem['h3FD9]=8'h00; mem['h3FDA]=8'h00; mem['h3FDB]=8'h00;
    mem['h3FDC]=8'h00; mem['h3FDD]=8'h00; mem['h3FDE]=8'h00; mem['h3FDF]=8'h00;
    mem['h3FE0]=8'h00; mem['h3FE1]=8'h00; mem['h3FE2]=8'h00; mem['h3FE3]=8'h00;
    mem['h3FE4]=8'h00; mem['h3FE5]=8'h00; mem['h3FE6]=8'h00; mem['h3FE7]=8'h00;
    mem['h3FE8]=8'h00; mem['h3FE9]=8'h00; mem['h3FEA]=8'h00; mem['h3FEB]=8'h00;
    mem['h3FEC]=8'h00; mem['h3FED]=8'h00; mem['h3FEE]=8'h00; mem['h3FEF]=8'h00;
    mem['h3FF0]=8'h00; mem['h3FF1]=8'h00; mem['h3FF2]=8'h00; mem['h3FF3]=8'h00;
    mem['h3FF4]=8'h00; mem['h3FF5]=8'h00; mem['h3FF6]=8'h00; mem['h3FF7]=8'h00;
    mem['h3FF8]=8'h00; mem['h3FF9]=8'h00; mem['h3FFA]=8'h00; mem['h3FFB]=8'h00;
    mem['h3FFC]=8'h00; mem['h3FFD]=8'h00; mem['h3FFE]=8'h00; mem['h3FFF]=8'h00;
    mem['h4000]=8'h00; mem['h4001]=8'h00; mem['h4002]=8'h00; mem['h4003]=8'h00;
    mem['h4004]=8'h00; mem['h4005]=8'h00; mem['h4006]=8'h00; mem['h4007]=8'h00;
    mem['h4008]=8'h00; mem['h4009]=8'h00; mem['h400A]=8'h00; mem['h400B]=8'h00;
    mem['h400C]=8'h00; mem['h400D]=8'h00; mem['h400E]=8'h00; mem['h400F]=8'h00;
    mem['h4010]=8'h00; mem['h4011]=8'h00; mem['h4012]=8'h00; mem['h4013]=8'h00;
    mem['h4014]=8'h00; mem['h4015]=8'h00; mem['h4016]=8'h00; mem['h4017]=8'h00;
    mem['h4018]=8'h00; mem['h4019]=8'h00; mem['h401A]=8'h00; mem['h401B]=8'h00;
    mem['h401C]=8'h00; mem['h401D]=8'h00; mem['h401E]=8'h00; mem['h401F]=8'h00;
    mem['h4020]=8'h00; mem['h4021]=8'h00; mem['h4022]=8'h00; mem['h4023]=8'h00;
    mem['h4024]=8'h00; mem['h4025]=8'h00; mem['h4026]=8'h00; mem['h4027]=8'h00;
    mem['h4028]=8'h00; mem['h4029]=8'h00; mem['h402A]=8'h00; mem['h402B]=8'h00;
    mem['h402C]=8'h00; mem['h402D]=8'h00; mem['h402E]=8'h00; mem['h402F]=8'h00;
    mem['h4030]=8'h00; mem['h4031]=8'h00; mem['h4032]=8'h00; mem['h4033]=8'h00;
    mem['h4034]=8'h00; mem['h4035]=8'h00; mem['h4036]=8'h00; mem['h4037]=8'h00;
    mem['h4038]=8'h00; mem['h4039]=8'h00; mem['h403A]=8'h00; mem['h403B]=8'h00;
    mem['h403C]=8'h00; mem['h403D]=8'h00; mem['h403E]=8'h00; mem['h403F]=8'h00;
    mem['h4040]=8'h00; mem['h4041]=8'h00; mem['h4042]=8'h00; mem['h4043]=8'h00;
    mem['h4044]=8'h00; mem['h4045]=8'h00; mem['h4046]=8'h00; mem['h4047]=8'h00;
    mem['h4048]=8'h00; mem['h4049]=8'h00; mem['h404A]=8'h00; mem['h404B]=8'h00;
    mem['h404C]=8'h00; mem['h404D]=8'h00; mem['h404E]=8'h00; mem['h404F]=8'h00;
    mem['h4050]=8'h00; mem['h4051]=8'h00; mem['h4052]=8'h00; mem['h4053]=8'h00;
    mem['h4054]=8'h00; mem['h4055]=8'h00; mem['h4056]=8'h00; mem['h4057]=8'h00;
    mem['h4058]=8'h00; mem['h4059]=8'h00; mem['h405A]=8'h00; mem['h405B]=8'h00;
    mem['h405C]=8'h00; mem['h405D]=8'h00; mem['h405E]=8'h00; mem['h405F]=8'h00;
    mem['h4060]=8'h00; mem['h4061]=8'h00; mem['h4062]=8'h00; mem['h4063]=8'h00;
    mem['h4064]=8'h00; mem['h4065]=8'h00; mem['h4066]=8'h00; mem['h4067]=8'h00;
    mem['h4068]=8'h00; mem['h4069]=8'h00; mem['h406A]=8'h00; mem['h406B]=8'h00;
    mem['h406C]=8'h00; mem['h406D]=8'h00; mem['h406E]=8'h00; mem['h406F]=8'h00;
    mem['h4070]=8'h00; mem['h4071]=8'h00; mem['h4072]=8'h00; mem['h4073]=8'h00;
    mem['h4074]=8'h00; mem['h4075]=8'h00; mem['h4076]=8'h00; mem['h4077]=8'h00;
    mem['h4078]=8'h00; mem['h4079]=8'h00; mem['h407A]=8'h00; mem['h407B]=8'h00;
    mem['h407C]=8'h00; mem['h407D]=8'h00; mem['h407E]=8'h00; mem['h407F]=8'h00;
    mem['h4080]=8'h00; mem['h4081]=8'h00; mem['h4082]=8'h00; mem['h4083]=8'h00;
    mem['h4084]=8'h00; mem['h4085]=8'h00; mem['h4086]=8'h00; mem['h4087]=8'h00;
    mem['h4088]=8'h00; mem['h4089]=8'h00; mem['h408A]=8'h00; mem['h408B]=8'h00;
    mem['h408C]=8'h00; mem['h408D]=8'h00; mem['h408E]=8'h00; mem['h408F]=8'h00;
    mem['h4090]=8'h00; mem['h4091]=8'h00; mem['h4092]=8'h00; mem['h4093]=8'h00;
    mem['h4094]=8'h00; mem['h4095]=8'h00; mem['h4096]=8'h00; mem['h4097]=8'h00;
    mem['h4098]=8'h00; mem['h4099]=8'h00; mem['h409A]=8'h00; mem['h409B]=8'h00;
    mem['h409C]=8'h00; mem['h409D]=8'h00; mem['h409E]=8'h00; mem['h409F]=8'h00;
    mem['h40A0]=8'h00; mem['h40A1]=8'h00; mem['h40A2]=8'h00; mem['h40A3]=8'h00;
    mem['h40A4]=8'h00; mem['h40A5]=8'h00; mem['h40A6]=8'h00; mem['h40A7]=8'h00;
    mem['h40A8]=8'h00; mem['h40A9]=8'h00; mem['h40AA]=8'h00; mem['h40AB]=8'h00;
    mem['h40AC]=8'h00; mem['h40AD]=8'h00; mem['h40AE]=8'h00; mem['h40AF]=8'h00;
    mem['h40B0]=8'h00; mem['h40B1]=8'h00; mem['h40B2]=8'h00; mem['h40B3]=8'h00;
    mem['h40B4]=8'h00; mem['h40B5]=8'h00; mem['h40B6]=8'h00; mem['h40B7]=8'h00;
    mem['h40B8]=8'h00; mem['h40B9]=8'h00; mem['h40BA]=8'h00; mem['h40BB]=8'h00;
    mem['h40BC]=8'h00; mem['h40BD]=8'h00; mem['h40BE]=8'h00; mem['h40BF]=8'h00;
    mem['h40C0]=8'h00; mem['h40C1]=8'h00; mem['h40C2]=8'h00; mem['h40C3]=8'h00;
    mem['h40C4]=8'h00; mem['h40C5]=8'h00; mem['h40C6]=8'h00; mem['h40C7]=8'h00;
    mem['h40C8]=8'h00; mem['h40C9]=8'h00; mem['h40CA]=8'h00; mem['h40CB]=8'h00;
    mem['h40CC]=8'h00; mem['h40CD]=8'h00; mem['h40CE]=8'h00; mem['h40CF]=8'h00;
    mem['h40D0]=8'h00; mem['h40D1]=8'h00; mem['h40D2]=8'h00; mem['h40D3]=8'h00;
    mem['h40D4]=8'h00; mem['h40D5]=8'h00; mem['h40D6]=8'h00; mem['h40D7]=8'h00;
    mem['h40D8]=8'h00; mem['h40D9]=8'h00; mem['h40DA]=8'h00; mem['h40DB]=8'h00;
    mem['h40DC]=8'h00; mem['h40DD]=8'h00; mem['h40DE]=8'h00; mem['h40DF]=8'h00;
    mem['h40E0]=8'h00; mem['h40E1]=8'h00; mem['h40E2]=8'h00; mem['h40E3]=8'h00;
    mem['h40E4]=8'h00; mem['h40E5]=8'h00; mem['h40E6]=8'h00; mem['h40E7]=8'h00;
    mem['h40E8]=8'h00; mem['h40E9]=8'h00; mem['h40EA]=8'h00; mem['h40EB]=8'h00;
    mem['h40EC]=8'h00; mem['h40ED]=8'h00; mem['h40EE]=8'h00; mem['h40EF]=8'h00;
    mem['h40F0]=8'h00; mem['h40F1]=8'h00; mem['h40F2]=8'h00; mem['h40F3]=8'h00;
    mem['h40F4]=8'h00; mem['h40F5]=8'h00; mem['h40F6]=8'h00; mem['h40F7]=8'h00;
    mem['h40F8]=8'h00; mem['h40F9]=8'h00; mem['h40FA]=8'h00; mem['h40FB]=8'h00;
    mem['h40FC]=8'h00; mem['h40FD]=8'h00; mem['h40FE]=8'h00; mem['h40FF]=8'h00;
    mem['h4100]=8'h00; mem['h4101]=8'h00; mem['h4102]=8'h00; mem['h4103]=8'h00;
    mem['h4104]=8'h00; mem['h4105]=8'h00; mem['h4106]=8'h00; mem['h4107]=8'h00;
    mem['h4108]=8'h00; mem['h4109]=8'h00; mem['h410A]=8'h00; mem['h410B]=8'h00;
    mem['h410C]=8'h00; mem['h410D]=8'h00; mem['h410E]=8'h00; mem['h410F]=8'h00;
    mem['h4110]=8'h00; mem['h4111]=8'h00; mem['h4112]=8'h00; mem['h4113]=8'h00;
    mem['h4114]=8'h00; mem['h4115]=8'h00; mem['h4116]=8'h00; mem['h4117]=8'h00;
    mem['h4118]=8'h00; mem['h4119]=8'h00; mem['h411A]=8'h00; mem['h411B]=8'h00;
    mem['h411C]=8'h00; mem['h411D]=8'h00; mem['h411E]=8'h00; mem['h411F]=8'h00;
    mem['h4120]=8'h00; mem['h4121]=8'h00; mem['h4122]=8'h00; mem['h4123]=8'h00;
    mem['h4124]=8'h00; mem['h4125]=8'h00; mem['h4126]=8'h00; mem['h4127]=8'h00;
    mem['h4128]=8'h00; mem['h4129]=8'h00; mem['h412A]=8'h00; mem['h412B]=8'h00;
    mem['h412C]=8'h00; mem['h412D]=8'h00; mem['h412E]=8'h00; mem['h412F]=8'h00;
    mem['h4130]=8'h00; mem['h4131]=8'h00; mem['h4132]=8'h00; mem['h4133]=8'h00;
    mem['h4134]=8'h00; mem['h4135]=8'h00; mem['h4136]=8'h00; mem['h4137]=8'h00;
    mem['h4138]=8'h00; mem['h4139]=8'h00; mem['h413A]=8'h00; mem['h413B]=8'h00;
    mem['h413C]=8'h00; mem['h413D]=8'h00; mem['h413E]=8'h00; mem['h413F]=8'h00;
    mem['h4140]=8'h00; mem['h4141]=8'h00; mem['h4142]=8'h00; mem['h4143]=8'h00;
    mem['h4144]=8'h00; mem['h4145]=8'h00; mem['h4146]=8'h00; mem['h4147]=8'h00;
    mem['h4148]=8'h00; mem['h4149]=8'h00; mem['h414A]=8'h00; mem['h414B]=8'h00;
    mem['h414C]=8'h00; mem['h414D]=8'h00; mem['h414E]=8'h00; mem['h414F]=8'h00;
    mem['h4150]=8'h00; mem['h4151]=8'h00; mem['h4152]=8'h00; mem['h4153]=8'h00;
    mem['h4154]=8'h00; mem['h4155]=8'h00; mem['h4156]=8'h00; mem['h4157]=8'h00;
    mem['h4158]=8'h00; mem['h4159]=8'h00; mem['h415A]=8'h00; mem['h415B]=8'h00;
    mem['h415C]=8'h00; mem['h415D]=8'h00; mem['h415E]=8'h00; mem['h415F]=8'h00;
    mem['h4160]=8'h00; mem['h4161]=8'h00; mem['h4162]=8'h00; mem['h4163]=8'h00;
    mem['h4164]=8'h00; mem['h4165]=8'h00; mem['h4166]=8'h00; mem['h4167]=8'h00;
    mem['h4168]=8'h00; mem['h4169]=8'h00; mem['h416A]=8'h00; mem['h416B]=8'h00;
    mem['h416C]=8'h00; mem['h416D]=8'h00; mem['h416E]=8'h00; mem['h416F]=8'h00;
    mem['h4170]=8'h00; mem['h4171]=8'h00; mem['h4172]=8'h00; mem['h4173]=8'h00;
    mem['h4174]=8'h00; mem['h4175]=8'h00; mem['h4176]=8'h00; mem['h4177]=8'h00;
    mem['h4178]=8'h00; mem['h4179]=8'h00; mem['h417A]=8'h00; mem['h417B]=8'h00;
    mem['h417C]=8'h00; mem['h417D]=8'h00; mem['h417E]=8'h00; mem['h417F]=8'h00;
    mem['h4180]=8'h00; mem['h4181]=8'h00; mem['h4182]=8'h00; mem['h4183]=8'h00;
    mem['h4184]=8'h00; mem['h4185]=8'h00; mem['h4186]=8'h00; mem['h4187]=8'h00;
    mem['h4188]=8'h00; mem['h4189]=8'h00; mem['h418A]=8'h00; mem['h418B]=8'h00;
    mem['h418C]=8'h00; mem['h418D]=8'h00; mem['h418E]=8'h00; mem['h418F]=8'h00;
    mem['h4190]=8'h00; mem['h4191]=8'h00; mem['h4192]=8'h00; mem['h4193]=8'h00;
    mem['h4194]=8'h00; mem['h4195]=8'h00; mem['h4196]=8'h00; mem['h4197]=8'h00;
    mem['h4198]=8'h00; mem['h4199]=8'h00; mem['h419A]=8'h00; mem['h419B]=8'h00;
    mem['h419C]=8'h00; mem['h419D]=8'h00; mem['h419E]=8'h00; mem['h419F]=8'h00;
    mem['h41A0]=8'h00; mem['h41A1]=8'h00; mem['h41A2]=8'h00; mem['h41A3]=8'h00;
    mem['h41A4]=8'h00; mem['h41A5]=8'h00; mem['h41A6]=8'h00; mem['h41A7]=8'h00;
    mem['h41A8]=8'h00; mem['h41A9]=8'h00; mem['h41AA]=8'h00; mem['h41AB]=8'h00;
    mem['h41AC]=8'h00; mem['h41AD]=8'h00; mem['h41AE]=8'h00; mem['h41AF]=8'h00;
    mem['h41B0]=8'h00; mem['h41B1]=8'h00; mem['h41B2]=8'h00; mem['h41B3]=8'h00;
    mem['h41B4]=8'h00; mem['h41B5]=8'h00; mem['h41B6]=8'h00; mem['h41B7]=8'h00;
    mem['h41B8]=8'h00; mem['h41B9]=8'h00; mem['h41BA]=8'h00; mem['h41BB]=8'h00;
    mem['h41BC]=8'h00; mem['h41BD]=8'h00; mem['h41BE]=8'h00; mem['h41BF]=8'h00;
    mem['h41C0]=8'h00; mem['h41C1]=8'h00; mem['h41C2]=8'h00; mem['h41C3]=8'h00;
    mem['h41C4]=8'h00; mem['h41C5]=8'h00; mem['h41C6]=8'h00; mem['h41C7]=8'h00;
    mem['h41C8]=8'h00; mem['h41C9]=8'h00; mem['h41CA]=8'h00; mem['h41CB]=8'h00;
    mem['h41CC]=8'h00; mem['h41CD]=8'h00; mem['h41CE]=8'h00; mem['h41CF]=8'h00;
    mem['h41D0]=8'h00; mem['h41D1]=8'h00; mem['h41D2]=8'h00; mem['h41D3]=8'h00;
    mem['h41D4]=8'h00; mem['h41D5]=8'h00; mem['h41D6]=8'h00; mem['h41D7]=8'h00;
    mem['h41D8]=8'h00; mem['h41D9]=8'h00; mem['h41DA]=8'h00; mem['h41DB]=8'h00;
    mem['h41DC]=8'h00; mem['h41DD]=8'h00; mem['h41DE]=8'h00; mem['h41DF]=8'h00;
    mem['h41E0]=8'h00; mem['h41E1]=8'h00; mem['h41E2]=8'h00; mem['h41E3]=8'h00;
    mem['h41E4]=8'h00; mem['h41E5]=8'h00; mem['h41E6]=8'h00; mem['h41E7]=8'h00;
    mem['h41E8]=8'h00; mem['h41E9]=8'h00; mem['h41EA]=8'h00; mem['h41EB]=8'h00;
    mem['h41EC]=8'h00; mem['h41ED]=8'h00; mem['h41EE]=8'h00; mem['h41EF]=8'h00;
    mem['h41F0]=8'h00; mem['h41F1]=8'h00; mem['h41F2]=8'h00; mem['h41F3]=8'h00;
    mem['h41F4]=8'h00; mem['h41F5]=8'h00; mem['h41F6]=8'h00; mem['h41F7]=8'h00;
    mem['h41F8]=8'h00; mem['h41F9]=8'h00; mem['h41FA]=8'h00; mem['h41FB]=8'h00;
    mem['h41FC]=8'h00; mem['h41FD]=8'h00; mem['h41FE]=8'h00; mem['h41FF]=8'h00;
    mem['h4200]=8'h00; mem['h4201]=8'h00; mem['h4202]=8'h00; mem['h4203]=8'h00;
    mem['h4204]=8'h00; mem['h4205]=8'h00; mem['h4206]=8'h00; mem['h4207]=8'h00;
    mem['h4208]=8'h00; mem['h4209]=8'h00; mem['h420A]=8'h00; mem['h420B]=8'h00;
    mem['h420C]=8'h00; mem['h420D]=8'h00; mem['h420E]=8'h00; mem['h420F]=8'h00;
    mem['h4210]=8'h00; mem['h4211]=8'h00; mem['h4212]=8'h00; mem['h4213]=8'h00;
    mem['h4214]=8'h00; mem['h4215]=8'h00; mem['h4216]=8'h00; mem['h4217]=8'h00;
    mem['h4218]=8'h00; mem['h4219]=8'h00; mem['h421A]=8'h00; mem['h421B]=8'h00;
    mem['h421C]=8'h00; mem['h421D]=8'h00; mem['h421E]=8'h00; mem['h421F]=8'h00;
    mem['h4220]=8'h00; mem['h4221]=8'h00; mem['h4222]=8'h00; mem['h4223]=8'h00;
    mem['h4224]=8'h00; mem['h4225]=8'h00; mem['h4226]=8'h00; mem['h4227]=8'h00;
    mem['h4228]=8'h00; mem['h4229]=8'h00; mem['h422A]=8'h00; mem['h422B]=8'h00;
    mem['h422C]=8'h00; mem['h422D]=8'h00; mem['h422E]=8'h00; mem['h422F]=8'h00;
    mem['h4230]=8'h00; mem['h4231]=8'h00; mem['h4232]=8'h00; mem['h4233]=8'h00;
    mem['h4234]=8'h00; mem['h4235]=8'h00; mem['h4236]=8'h00; mem['h4237]=8'h00;
    mem['h4238]=8'h00; mem['h4239]=8'h00; mem['h423A]=8'h00; mem['h423B]=8'h00;
    mem['h423C]=8'h00; mem['h423D]=8'h00; mem['h423E]=8'h00; mem['h423F]=8'h00;
    mem['h4240]=8'h00; mem['h4241]=8'h00; mem['h4242]=8'h00; mem['h4243]=8'h00;
    mem['h4244]=8'h00; mem['h4245]=8'h00; mem['h4246]=8'h00; mem['h4247]=8'h00;
    mem['h4248]=8'h00; mem['h4249]=8'h00; mem['h424A]=8'h00; mem['h424B]=8'h00;
    mem['h424C]=8'h00; mem['h424D]=8'h00; mem['h424E]=8'h00; mem['h424F]=8'h00;
    mem['h4250]=8'h00; mem['h4251]=8'h00; mem['h4252]=8'h00; mem['h4253]=8'h00;
    mem['h4254]=8'h00; mem['h4255]=8'h00; mem['h4256]=8'h00; mem['h4257]=8'h00;
    mem['h4258]=8'h00; mem['h4259]=8'h00; mem['h425A]=8'h00; mem['h425B]=8'h00;
    mem['h425C]=8'h00; mem['h425D]=8'h00; mem['h425E]=8'h00; mem['h425F]=8'h00;
    mem['h4260]=8'h00; mem['h4261]=8'h00; mem['h4262]=8'h00; mem['h4263]=8'h00;
    mem['h4264]=8'h00; mem['h4265]=8'h00; mem['h4266]=8'h00; mem['h4267]=8'h00;
    mem['h4268]=8'h00; mem['h4269]=8'h00; mem['h426A]=8'h00; mem['h426B]=8'h00;
    mem['h426C]=8'h00; mem['h426D]=8'h00; mem['h426E]=8'h00; mem['h426F]=8'h00;
    mem['h4270]=8'h00; mem['h4271]=8'h00; mem['h4272]=8'h00; mem['h4273]=8'h00;
    mem['h4274]=8'h00; mem['h4275]=8'h00; mem['h4276]=8'h00; mem['h4277]=8'h00;
    mem['h4278]=8'h00; mem['h4279]=8'h00; mem['h427A]=8'h00; mem['h427B]=8'h00;
    mem['h427C]=8'h00; mem['h427D]=8'h00; mem['h427E]=8'h00; mem['h427F]=8'h00;
    mem['h4280]=8'h00; mem['h4281]=8'h00; mem['h4282]=8'h00; mem['h4283]=8'h00;
    mem['h4284]=8'h00; mem['h4285]=8'h00; mem['h4286]=8'h00; mem['h4287]=8'h00;
    mem['h4288]=8'h00; mem['h4289]=8'h00; mem['h428A]=8'h00; mem['h428B]=8'h00;
    mem['h428C]=8'h00; mem['h428D]=8'h00; mem['h428E]=8'h00; mem['h428F]=8'h00;
    mem['h4290]=8'h00; mem['h4291]=8'h00; mem['h4292]=8'h00; mem['h4293]=8'h00;
    mem['h4294]=8'h00; mem['h4295]=8'h00; mem['h4296]=8'h00; mem['h4297]=8'h00;
    mem['h4298]=8'h00; mem['h4299]=8'h00; mem['h429A]=8'h00; mem['h429B]=8'h00;
    mem['h429C]=8'h00; mem['h429D]=8'h00; mem['h429E]=8'h00; mem['h429F]=8'h00;
    mem['h42A0]=8'h00; mem['h42A1]=8'h00; mem['h42A2]=8'h00; mem['h42A3]=8'h00;
    mem['h42A4]=8'h00; mem['h42A5]=8'h00; mem['h42A6]=8'h00; mem['h42A7]=8'h00;
    mem['h42A8]=8'h00; mem['h42A9]=8'h00; mem['h42AA]=8'h00; mem['h42AB]=8'h00;
    mem['h42AC]=8'h00; mem['h42AD]=8'h00; mem['h42AE]=8'h00; mem['h42AF]=8'h00;
    mem['h42B0]=8'h00; mem['h42B1]=8'h00; mem['h42B2]=8'h00; mem['h42B3]=8'h00;
    mem['h42B4]=8'h00; mem['h42B5]=8'h00; mem['h42B6]=8'h00; mem['h42B7]=8'h00;
    mem['h42B8]=8'h00; mem['h42B9]=8'h00; mem['h42BA]=8'h00; mem['h42BB]=8'h00;
    mem['h42BC]=8'h00; mem['h42BD]=8'h00; mem['h42BE]=8'h00; mem['h42BF]=8'h00;
    mem['h42C0]=8'h00; mem['h42C1]=8'h00; mem['h42C2]=8'h00; mem['h42C3]=8'h00;
    mem['h42C4]=8'h00; mem['h42C5]=8'h00; mem['h42C6]=8'h00; mem['h42C7]=8'h00;
    mem['h42C8]=8'h00; mem['h42C9]=8'h00; mem['h42CA]=8'h00; mem['h42CB]=8'h00;
    mem['h42CC]=8'h00; mem['h42CD]=8'h00; mem['h42CE]=8'h00; mem['h42CF]=8'h00;
    mem['h42D0]=8'h00; mem['h42D1]=8'h00; mem['h42D2]=8'h00; mem['h42D3]=8'h00;
    mem['h42D4]=8'h00; mem['h42D5]=8'h00; mem['h42D6]=8'h00; mem['h42D7]=8'h00;
    mem['h42D8]=8'h00; mem['h42D9]=8'h00; mem['h42DA]=8'h00; mem['h42DB]=8'h00;
    mem['h42DC]=8'h00; mem['h42DD]=8'h00; mem['h42DE]=8'h00; mem['h42DF]=8'h00;
    mem['h42E0]=8'h00; mem['h42E1]=8'h00; mem['h42E2]=8'h00; mem['h42E3]=8'h00;
    mem['h42E4]=8'h00; mem['h42E5]=8'h00; mem['h42E6]=8'h00; mem['h42E7]=8'h00;
    mem['h42E8]=8'h00; mem['h42E9]=8'h00; mem['h42EA]=8'h00; mem['h42EB]=8'h00;
    mem['h42EC]=8'h00; mem['h42ED]=8'h00; mem['h42EE]=8'h00; mem['h42EF]=8'h00;
    mem['h42F0]=8'h00; mem['h42F1]=8'h00; mem['h42F2]=8'h00; mem['h42F3]=8'h00;
    mem['h42F4]=8'h00; mem['h42F5]=8'h00; mem['h42F6]=8'h00; mem['h42F7]=8'h00;
    mem['h42F8]=8'h00; mem['h42F9]=8'h00; mem['h42FA]=8'h00; mem['h42FB]=8'h00;
    mem['h42FC]=8'h00; mem['h42FD]=8'h00; mem['h42FE]=8'h00; mem['h42FF]=8'h00;
    mem['h4300]=8'h00; mem['h4301]=8'h00; mem['h4302]=8'h00; mem['h4303]=8'h00;
    mem['h4304]=8'h00; mem['h4305]=8'h00; mem['h4306]=8'h00; mem['h4307]=8'h00;
    mem['h4308]=8'h00; mem['h4309]=8'h00; mem['h430A]=8'h00; mem['h430B]=8'h00;
    mem['h430C]=8'h00; mem['h430D]=8'h00; mem['h430E]=8'h00; mem['h430F]=8'h00;
    mem['h4310]=8'h00; mem['h4311]=8'h00; mem['h4312]=8'h00; mem['h4313]=8'h00;
    mem['h4314]=8'h00; mem['h4315]=8'h00; mem['h4316]=8'h00; mem['h4317]=8'h00;
    mem['h4318]=8'h00; mem['h4319]=8'h00; mem['h431A]=8'h00; mem['h431B]=8'h00;
    mem['h431C]=8'h00; mem['h431D]=8'h00; mem['h431E]=8'h00; mem['h431F]=8'h00;
    mem['h4320]=8'h00; mem['h4321]=8'h00; mem['h4322]=8'h00; mem['h4323]=8'h00;
    mem['h4324]=8'h00; mem['h4325]=8'h00; mem['h4326]=8'h00; mem['h4327]=8'h00;
    mem['h4328]=8'h00; mem['h4329]=8'h00; mem['h432A]=8'h00; mem['h432B]=8'h00;
    mem['h432C]=8'h00; mem['h432D]=8'h00; mem['h432E]=8'h00; mem['h432F]=8'h00;
    mem['h4330]=8'h00; mem['h4331]=8'h00; mem['h4332]=8'h00; mem['h4333]=8'h00;
    mem['h4334]=8'h00; mem['h4335]=8'h00; mem['h4336]=8'h00; mem['h4337]=8'h00;
    mem['h4338]=8'h00; mem['h4339]=8'h00; mem['h433A]=8'h00; mem['h433B]=8'h00;
    mem['h433C]=8'h00; mem['h433D]=8'h00; mem['h433E]=8'h00; mem['h433F]=8'h00;
    mem['h4340]=8'h00; mem['h4341]=8'h00; mem['h4342]=8'h00; mem['h4343]=8'h00;
    mem['h4344]=8'h00; mem['h4345]=8'h00; mem['h4346]=8'h00; mem['h4347]=8'h00;
    mem['h4348]=8'h00; mem['h4349]=8'h00; mem['h434A]=8'h00; mem['h434B]=8'h00;
    mem['h434C]=8'h00; mem['h434D]=8'h00; mem['h434E]=8'h00; mem['h434F]=8'h00;
    mem['h4350]=8'h00; mem['h4351]=8'h00; mem['h4352]=8'h00; mem['h4353]=8'h00;
    mem['h4354]=8'h00; mem['h4355]=8'h00; mem['h4356]=8'h00; mem['h4357]=8'h00;
    mem['h4358]=8'h00; mem['h4359]=8'h00; mem['h435A]=8'h00; mem['h435B]=8'h00;
    mem['h435C]=8'h00; mem['h435D]=8'h00; mem['h435E]=8'h00; mem['h435F]=8'h00;
    mem['h4360]=8'h00; mem['h4361]=8'h00; mem['h4362]=8'h00; mem['h4363]=8'h00;
    mem['h4364]=8'h00; mem['h4365]=8'h00; mem['h4366]=8'h00; mem['h4367]=8'h00;
    mem['h4368]=8'h00; mem['h4369]=8'h00; mem['h436A]=8'h00; mem['h436B]=8'h00;
    mem['h436C]=8'h00; mem['h436D]=8'h00; mem['h436E]=8'h00; mem['h436F]=8'h00;
    mem['h4370]=8'h00; mem['h4371]=8'h00; mem['h4372]=8'h00; mem['h4373]=8'h00;
    mem['h4374]=8'h00; mem['h4375]=8'h00; mem['h4376]=8'h00; mem['h4377]=8'h00;
    mem['h4378]=8'h00; mem['h4379]=8'h00; mem['h437A]=8'h00; mem['h437B]=8'h00;
    mem['h437C]=8'h00; mem['h437D]=8'h00; mem['h437E]=8'h00; mem['h437F]=8'h00;
    mem['h4380]=8'h00; mem['h4381]=8'h00; mem['h4382]=8'h00; mem['h4383]=8'h00;
    mem['h4384]=8'h00; mem['h4385]=8'h00; mem['h4386]=8'h00; mem['h4387]=8'h00;
    mem['h4388]=8'h00; mem['h4389]=8'h00; mem['h438A]=8'h00; mem['h438B]=8'h00;
    mem['h438C]=8'h00; mem['h438D]=8'h00; mem['h438E]=8'h00; mem['h438F]=8'h00;
    mem['h4390]=8'h00; mem['h4391]=8'h00; mem['h4392]=8'h00; mem['h4393]=8'h00;
    mem['h4394]=8'h00; mem['h4395]=8'h00; mem['h4396]=8'h00; mem['h4397]=8'h00;
    mem['h4398]=8'h00; mem['h4399]=8'h00; mem['h439A]=8'h00; mem['h439B]=8'h00;
    mem['h439C]=8'h00; mem['h439D]=8'h00; mem['h439E]=8'h00; mem['h439F]=8'h00;
    mem['h43A0]=8'h00; mem['h43A1]=8'h00; mem['h43A2]=8'h00; mem['h43A3]=8'h00;
    mem['h43A4]=8'h00; mem['h43A5]=8'h00; mem['h43A6]=8'h00; mem['h43A7]=8'h00;
    mem['h43A8]=8'h00; mem['h43A9]=8'h00; mem['h43AA]=8'h00; mem['h43AB]=8'h00;
    mem['h43AC]=8'h00; mem['h43AD]=8'h00; mem['h43AE]=8'h00; mem['h43AF]=8'h00;
    mem['h43B0]=8'h00; mem['h43B1]=8'h00; mem['h43B2]=8'h00; mem['h43B3]=8'h00;
    mem['h43B4]=8'h00; mem['h43B5]=8'h00; mem['h43B6]=8'h00; mem['h43B7]=8'h00;
    mem['h43B8]=8'h00; mem['h43B9]=8'h00; mem['h43BA]=8'h00; mem['h43BB]=8'h00;
    mem['h43BC]=8'h00; mem['h43BD]=8'h00; mem['h43BE]=8'h00; mem['h43BF]=8'h00;
    mem['h43C0]=8'h00; mem['h43C1]=8'h00; mem['h43C2]=8'h00; mem['h43C3]=8'h00;
    mem['h43C4]=8'h00; mem['h43C5]=8'h00; mem['h43C6]=8'h00; mem['h43C7]=8'h00;
    mem['h43C8]=8'h00; mem['h43C9]=8'h00; mem['h43CA]=8'h00; mem['h43CB]=8'h00;
    mem['h43CC]=8'h00; mem['h43CD]=8'h00; mem['h43CE]=8'h00; mem['h43CF]=8'h00;
    mem['h43D0]=8'h00; mem['h43D1]=8'h00; mem['h43D2]=8'h00; mem['h43D3]=8'h00;
    mem['h43D4]=8'h00; mem['h43D5]=8'h00; mem['h43D6]=8'h00; mem['h43D7]=8'h00;
    mem['h43D8]=8'h00; mem['h43D9]=8'h00; mem['h43DA]=8'h00; mem['h43DB]=8'h00;
    mem['h43DC]=8'h00; mem['h43DD]=8'h00; mem['h43DE]=8'h00; mem['h43DF]=8'h00;
    mem['h43E0]=8'h00; mem['h43E1]=8'h00; mem['h43E2]=8'h00; mem['h43E3]=8'h00;
    mem['h43E4]=8'h00; mem['h43E5]=8'h00; mem['h43E6]=8'h00; mem['h43E7]=8'h00;
    mem['h43E8]=8'h00; mem['h43E9]=8'h00; mem['h43EA]=8'h00; mem['h43EB]=8'h00;
    mem['h43EC]=8'h00; mem['h43ED]=8'h00; mem['h43EE]=8'h00; mem['h43EF]=8'h00;
    mem['h43F0]=8'h00; mem['h43F1]=8'h00; mem['h43F2]=8'h00; mem['h43F3]=8'h00;
    mem['h43F4]=8'h00; mem['h43F5]=8'h00; mem['h43F6]=8'h00; mem['h43F7]=8'h00;
    mem['h43F8]=8'h00; mem['h43F9]=8'h00; mem['h43FA]=8'h00; mem['h43FB]=8'h00;
    mem['h43FC]=8'h00; mem['h43FD]=8'h00; mem['h43FE]=8'h00; mem['h43FF]=8'h00;
    mem['h4400]=8'h00; mem['h4401]=8'h00; mem['h4402]=8'h00; mem['h4403]=8'h00;
    mem['h4404]=8'h00; mem['h4405]=8'h00; mem['h4406]=8'h00; mem['h4407]=8'h00;
    mem['h4408]=8'h00; mem['h4409]=8'h00; mem['h440A]=8'h00; mem['h440B]=8'h00;
    mem['h440C]=8'h00; mem['h440D]=8'h00; mem['h440E]=8'h00; mem['h440F]=8'h00;
    mem['h4410]=8'h00; mem['h4411]=8'h00; mem['h4412]=8'h00; mem['h4413]=8'h00;
    mem['h4414]=8'h00; mem['h4415]=8'h00; mem['h4416]=8'h00; mem['h4417]=8'h00;
    mem['h4418]=8'h00; mem['h4419]=8'h00; mem['h441A]=8'h00; mem['h441B]=8'h00;
    mem['h441C]=8'h00; mem['h441D]=8'h00; mem['h441E]=8'h00; mem['h441F]=8'h00;
    mem['h4420]=8'h00; mem['h4421]=8'h00; mem['h4422]=8'h00; mem['h4423]=8'h00;
    mem['h4424]=8'h00; mem['h4425]=8'h00; mem['h4426]=8'h00; mem['h4427]=8'h00;
    mem['h4428]=8'h00; mem['h4429]=8'h00; mem['h442A]=8'h00; mem['h442B]=8'h00;
    mem['h442C]=8'h00; mem['h442D]=8'h00; mem['h442E]=8'h00; mem['h442F]=8'h00;
    mem['h4430]=8'h00; mem['h4431]=8'h00; mem['h4432]=8'h00; mem['h4433]=8'h00;
    mem['h4434]=8'h00; mem['h4435]=8'h00; mem['h4436]=8'h00; mem['h4437]=8'h00;
    mem['h4438]=8'h00; mem['h4439]=8'h00; mem['h443A]=8'h00; mem['h443B]=8'h00;
    mem['h443C]=8'h00; mem['h443D]=8'h00; mem['h443E]=8'h00; mem['h443F]=8'h00;
    mem['h4440]=8'h00; mem['h4441]=8'h00; mem['h4442]=8'h00; mem['h4443]=8'h00;
    mem['h4444]=8'h00; mem['h4445]=8'h00; mem['h4446]=8'h00; mem['h4447]=8'h00;
    mem['h4448]=8'h00; mem['h4449]=8'h00; mem['h444A]=8'h00; mem['h444B]=8'h00;
    mem['h444C]=8'h00; mem['h444D]=8'h00; mem['h444E]=8'h00; mem['h444F]=8'h00;
    mem['h4450]=8'h00; mem['h4451]=8'h00; mem['h4452]=8'h00; mem['h4453]=8'h00;
    mem['h4454]=8'h00; mem['h4455]=8'h00; mem['h4456]=8'h00; mem['h4457]=8'h00;
    mem['h4458]=8'h00; mem['h4459]=8'h00; mem['h445A]=8'h00; mem['h445B]=8'h00;
    mem['h445C]=8'h00; mem['h445D]=8'h00; mem['h445E]=8'h00; mem['h445F]=8'h00;
    mem['h4460]=8'h00; mem['h4461]=8'h00; mem['h4462]=8'h00; mem['h4463]=8'h00;
    mem['h4464]=8'h00; mem['h4465]=8'h00; mem['h4466]=8'h00; mem['h4467]=8'h00;
    mem['h4468]=8'h00; mem['h4469]=8'h00; mem['h446A]=8'h00; mem['h446B]=8'h00;
    mem['h446C]=8'h00; mem['h446D]=8'h00; mem['h446E]=8'h00; mem['h446F]=8'h00;
    mem['h4470]=8'h00; mem['h4471]=8'h00; mem['h4472]=8'h00; mem['h4473]=8'h00;
    mem['h4474]=8'h00; mem['h4475]=8'h00; mem['h4476]=8'h00; mem['h4477]=8'h00;
    mem['h4478]=8'h00; mem['h4479]=8'h00; mem['h447A]=8'h00; mem['h447B]=8'h00;
    mem['h447C]=8'h00; mem['h447D]=8'h00; mem['h447E]=8'h00; mem['h447F]=8'h00;
    mem['h4480]=8'h00; mem['h4481]=8'h00; mem['h4482]=8'h00; mem['h4483]=8'h00;
    mem['h4484]=8'h00; mem['h4485]=8'h00; mem['h4486]=8'h00; mem['h4487]=8'h00;
    mem['h4488]=8'h00; mem['h4489]=8'h00; mem['h448A]=8'h00; mem['h448B]=8'h00;
    mem['h448C]=8'h00; mem['h448D]=8'h00; mem['h448E]=8'h00; mem['h448F]=8'h00;
    mem['h4490]=8'h00; mem['h4491]=8'h00; mem['h4492]=8'h00; mem['h4493]=8'h00;
    mem['h4494]=8'h00; mem['h4495]=8'h00; mem['h4496]=8'h00; mem['h4497]=8'h00;
    mem['h4498]=8'h00; mem['h4499]=8'h00; mem['h449A]=8'h00; mem['h449B]=8'h00;
    mem['h449C]=8'h00; mem['h449D]=8'h00; mem['h449E]=8'h00; mem['h449F]=8'h00;
    mem['h44A0]=8'h00; mem['h44A1]=8'h00; mem['h44A2]=8'h00; mem['h44A3]=8'h00;
    mem['h44A4]=8'h00; mem['h44A5]=8'h00; mem['h44A6]=8'h00; mem['h44A7]=8'h00;
    mem['h44A8]=8'h00; mem['h44A9]=8'h00; mem['h44AA]=8'h00; mem['h44AB]=8'h00;
    mem['h44AC]=8'h00; mem['h44AD]=8'h00; mem['h44AE]=8'h00; mem['h44AF]=8'h00;
    mem['h44B0]=8'h00; mem['h44B1]=8'h00; mem['h44B2]=8'h00; mem['h44B3]=8'h00;
    mem['h44B4]=8'h00; mem['h44B5]=8'h00; mem['h44B6]=8'h00; mem['h44B7]=8'h00;
    mem['h44B8]=8'h00; mem['h44B9]=8'h00; mem['h44BA]=8'h00; mem['h44BB]=8'h00;
    mem['h44BC]=8'h00; mem['h44BD]=8'h00; mem['h44BE]=8'h00; mem['h44BF]=8'h00;
    mem['h44C0]=8'h00; mem['h44C1]=8'h00; mem['h44C2]=8'h00; mem['h44C3]=8'h00;
    mem['h44C4]=8'h00; mem['h44C5]=8'h00; mem['h44C6]=8'h00; mem['h44C7]=8'h00;
    mem['h44C8]=8'h00; mem['h44C9]=8'h00; mem['h44CA]=8'h00; mem['h44CB]=8'h00;
    mem['h44CC]=8'h00; mem['h44CD]=8'h00; mem['h44CE]=8'h00; mem['h44CF]=8'h00;
    mem['h44D0]=8'h00; mem['h44D1]=8'h00; mem['h44D2]=8'h00; mem['h44D3]=8'h00;
    mem['h44D4]=8'h00; mem['h44D5]=8'h00; mem['h44D6]=8'h00; mem['h44D7]=8'h00;
    mem['h44D8]=8'h00; mem['h44D9]=8'h00; mem['h44DA]=8'h00; mem['h44DB]=8'h00;
    mem['h44DC]=8'h00; mem['h44DD]=8'h00; mem['h44DE]=8'h00; mem['h44DF]=8'h00;
    mem['h44E0]=8'h00; mem['h44E1]=8'h00; mem['h44E2]=8'h00; mem['h44E3]=8'h00;
    mem['h44E4]=8'h00; mem['h44E5]=8'h00; mem['h44E6]=8'h00; mem['h44E7]=8'h00;
    mem['h44E8]=8'h00; mem['h44E9]=8'h00; mem['h44EA]=8'h00; mem['h44EB]=8'h00;
    mem['h44EC]=8'h00; mem['h44ED]=8'h00; mem['h44EE]=8'h00; mem['h44EF]=8'h00;
    mem['h44F0]=8'h00; mem['h44F1]=8'h00; mem['h44F2]=8'h00; mem['h44F3]=8'h00;
    mem['h44F4]=8'h00; mem['h44F5]=8'h00; mem['h44F6]=8'h00; mem['h44F7]=8'h00;
    mem['h44F8]=8'h00; mem['h44F9]=8'h00; mem['h44FA]=8'h00; mem['h44FB]=8'h00;
    mem['h44FC]=8'h00; mem['h44FD]=8'h00; mem['h44FE]=8'h00; mem['h44FF]=8'h00;
    mem['h4500]=8'h00; mem['h4501]=8'h00; mem['h4502]=8'h00; mem['h4503]=8'h00;
    mem['h4504]=8'h00; mem['h4505]=8'h00; mem['h4506]=8'h00; mem['h4507]=8'h00;
    mem['h4508]=8'h00; mem['h4509]=8'h00; mem['h450A]=8'h00; mem['h450B]=8'h00;
    mem['h450C]=8'h00; mem['h450D]=8'h00; mem['h450E]=8'h00; mem['h450F]=8'h00;
    mem['h4510]=8'h00; mem['h4511]=8'h00; mem['h4512]=8'h00; mem['h4513]=8'h00;
    mem['h4514]=8'h00; mem['h4515]=8'h00; mem['h4516]=8'h00; mem['h4517]=8'h00;
    mem['h4518]=8'h00; mem['h4519]=8'h00; mem['h451A]=8'h00; mem['h451B]=8'h00;
    mem['h451C]=8'h00; mem['h451D]=8'h00; mem['h451E]=8'h00; mem['h451F]=8'h00;
    mem['h4520]=8'h00; mem['h4521]=8'h00; mem['h4522]=8'h00; mem['h4523]=8'h00;
    mem['h4524]=8'h00; mem['h4525]=8'h00; mem['h4526]=8'h00; mem['h4527]=8'h00;
    mem['h4528]=8'h00; mem['h4529]=8'h00; mem['h452A]=8'h00; mem['h452B]=8'h00;
    mem['h452C]=8'h00; mem['h452D]=8'h00; mem['h452E]=8'h00; mem['h452F]=8'h00;
    mem['h4530]=8'h00; mem['h4531]=8'h00; mem['h4532]=8'h00; mem['h4533]=8'h00;
    mem['h4534]=8'h00; mem['h4535]=8'h00; mem['h4536]=8'h00; mem['h4537]=8'h00;
    mem['h4538]=8'h00; mem['h4539]=8'h00; mem['h453A]=8'h00; mem['h453B]=8'h00;
    mem['h453C]=8'h00; mem['h453D]=8'h00; mem['h453E]=8'h00; mem['h453F]=8'h00;
    mem['h4540]=8'h00; mem['h4541]=8'h00; mem['h4542]=8'h00; mem['h4543]=8'h00;
    mem['h4544]=8'h00; mem['h4545]=8'h00; mem['h4546]=8'h00; mem['h4547]=8'h00;
    mem['h4548]=8'h00; mem['h4549]=8'h00; mem['h454A]=8'h00; mem['h454B]=8'h00;
    mem['h454C]=8'h00; mem['h454D]=8'h00; mem['h454E]=8'h00; mem['h454F]=8'h00;
    mem['h4550]=8'h00; mem['h4551]=8'h00; mem['h4552]=8'h00; mem['h4553]=8'h00;
    mem['h4554]=8'h00; mem['h4555]=8'h00; mem['h4556]=8'h00; mem['h4557]=8'h00;
    mem['h4558]=8'h00; mem['h4559]=8'h00; mem['h455A]=8'h00; mem['h455B]=8'h00;
    mem['h455C]=8'h00; mem['h455D]=8'h00; mem['h455E]=8'h00; mem['h455F]=8'h00;
    mem['h4560]=8'h00; mem['h4561]=8'h00; mem['h4562]=8'h00; mem['h4563]=8'h00;
    mem['h4564]=8'h00; mem['h4565]=8'h00; mem['h4566]=8'h00; mem['h4567]=8'h00;
    mem['h4568]=8'h00; mem['h4569]=8'h00; mem['h456A]=8'h00; mem['h456B]=8'h00;
    mem['h456C]=8'h00; mem['h456D]=8'h00; mem['h456E]=8'h00; mem['h456F]=8'h00;
    mem['h4570]=8'h00; mem['h4571]=8'h00; mem['h4572]=8'h00; mem['h4573]=8'h00;
    mem['h4574]=8'h00; mem['h4575]=8'h00; mem['h4576]=8'h00; mem['h4577]=8'h00;
    mem['h4578]=8'h00; mem['h4579]=8'h00; mem['h457A]=8'h00; mem['h457B]=8'h00;
    mem['h457C]=8'h00; mem['h457D]=8'h00; mem['h457E]=8'h00; mem['h457F]=8'h00;
    mem['h4580]=8'h00; mem['h4581]=8'h00; mem['h4582]=8'h00; mem['h4583]=8'h00;
    mem['h4584]=8'h00; mem['h4585]=8'h00; mem['h4586]=8'h00; mem['h4587]=8'h00;
    mem['h4588]=8'h00; mem['h4589]=8'h00; mem['h458A]=8'h00; mem['h458B]=8'h00;
    mem['h458C]=8'h00; mem['h458D]=8'h00; mem['h458E]=8'h00; mem['h458F]=8'h00;
    mem['h4590]=8'h00; mem['h4591]=8'h00; mem['h4592]=8'h00; mem['h4593]=8'h00;
    mem['h4594]=8'h00; mem['h4595]=8'h00; mem['h4596]=8'h00; mem['h4597]=8'h00;
    mem['h4598]=8'h00; mem['h4599]=8'h00; mem['h459A]=8'h00; mem['h459B]=8'h00;
    mem['h459C]=8'h00; mem['h459D]=8'h00; mem['h459E]=8'h00; mem['h459F]=8'h00;
    mem['h45A0]=8'h00; mem['h45A1]=8'h00; mem['h45A2]=8'h00; mem['h45A3]=8'h00;
    mem['h45A4]=8'h00; mem['h45A5]=8'h00; mem['h45A6]=8'h00; mem['h45A7]=8'h00;
    mem['h45A8]=8'h00; mem['h45A9]=8'h00; mem['h45AA]=8'h00; mem['h45AB]=8'h00;
    mem['h45AC]=8'h00; mem['h45AD]=8'h00; mem['h45AE]=8'h00; mem['h45AF]=8'h00;
    mem['h45B0]=8'h00; mem['h45B1]=8'h00; mem['h45B2]=8'h00; mem['h45B3]=8'h00;
    mem['h45B4]=8'h00; mem['h45B5]=8'h00; mem['h45B6]=8'h00; mem['h45B7]=8'h00;
    mem['h45B8]=8'h00; mem['h45B9]=8'h00; mem['h45BA]=8'h00; mem['h45BB]=8'h00;
    mem['h45BC]=8'h00; mem['h45BD]=8'h00; mem['h45BE]=8'h00; mem['h45BF]=8'h00;
    mem['h45C0]=8'h00; mem['h45C1]=8'h00; mem['h45C2]=8'h00; mem['h45C3]=8'h00;
    mem['h45C4]=8'h00; mem['h45C5]=8'h00; mem['h45C6]=8'h00; mem['h45C7]=8'h00;
    mem['h45C8]=8'h00; mem['h45C9]=8'h00; mem['h45CA]=8'h00; mem['h45CB]=8'h00;
    mem['h45CC]=8'h00; mem['h45CD]=8'h00; mem['h45CE]=8'h00; mem['h45CF]=8'h00;
    mem['h45D0]=8'h00; mem['h45D1]=8'h00; mem['h45D2]=8'h00; mem['h45D3]=8'h00;
    mem['h45D4]=8'h00; mem['h45D5]=8'h00; mem['h45D6]=8'h00; mem['h45D7]=8'h00;
    mem['h45D8]=8'h00; mem['h45D9]=8'h00; mem['h45DA]=8'h00; mem['h45DB]=8'h00;
    mem['h45DC]=8'h00; mem['h45DD]=8'h00; mem['h45DE]=8'h00; mem['h45DF]=8'h00;
    mem['h45E0]=8'h00; mem['h45E1]=8'h00; mem['h45E2]=8'h00; mem['h45E3]=8'h00;
    mem['h45E4]=8'h00; mem['h45E5]=8'h00; mem['h45E6]=8'h00; mem['h45E7]=8'h00;
    mem['h45E8]=8'h00; mem['h45E9]=8'h00; mem['h45EA]=8'h00; mem['h45EB]=8'h00;
    mem['h45EC]=8'h00; mem['h45ED]=8'h00; mem['h45EE]=8'h00; mem['h45EF]=8'h00;
    mem['h45F0]=8'h00; mem['h45F1]=8'h00; mem['h45F2]=8'h00; mem['h45F3]=8'h00;
    mem['h45F4]=8'h00; mem['h45F5]=8'h00; mem['h45F6]=8'h00; mem['h45F7]=8'h00;
    mem['h45F8]=8'h00; mem['h45F9]=8'h00; mem['h45FA]=8'h00; mem['h45FB]=8'h00;
    mem['h45FC]=8'h00; mem['h45FD]=8'h00; mem['h45FE]=8'h00; mem['h45FF]=8'h00;
    mem['h4600]=8'h00; mem['h4601]=8'h00; mem['h4602]=8'h00; mem['h4603]=8'h00;
    mem['h4604]=8'h00; mem['h4605]=8'h00; mem['h4606]=8'h00; mem['h4607]=8'h00;
    mem['h4608]=8'h00; mem['h4609]=8'h00; mem['h460A]=8'h00; mem['h460B]=8'h00;
    mem['h460C]=8'h00; mem['h460D]=8'h00; mem['h460E]=8'h00; mem['h460F]=8'h00;
    mem['h4610]=8'h00; mem['h4611]=8'h00; mem['h4612]=8'h00; mem['h4613]=8'h00;
    mem['h4614]=8'h00; mem['h4615]=8'h00; mem['h4616]=8'h00; mem['h4617]=8'h00;
    mem['h4618]=8'h00; mem['h4619]=8'h00; mem['h461A]=8'h00; mem['h461B]=8'h00;
    mem['h461C]=8'h00; mem['h461D]=8'h00; mem['h461E]=8'h00; mem['h461F]=8'h00;
    mem['h4620]=8'h00; mem['h4621]=8'h00; mem['h4622]=8'h00; mem['h4623]=8'h00;
    mem['h4624]=8'h00; mem['h4625]=8'h00; mem['h4626]=8'h00; mem['h4627]=8'h00;
    mem['h4628]=8'h00; mem['h4629]=8'h00; mem['h462A]=8'h00; mem['h462B]=8'h00;
    mem['h462C]=8'h00; mem['h462D]=8'h00; mem['h462E]=8'h00; mem['h462F]=8'h00;
    mem['h4630]=8'h00; mem['h4631]=8'h00; mem['h4632]=8'h00; mem['h4633]=8'h00;
    mem['h4634]=8'h00; mem['h4635]=8'h00; mem['h4636]=8'h00; mem['h4637]=8'h00;
    mem['h4638]=8'h00; mem['h4639]=8'h00; mem['h463A]=8'h00; mem['h463B]=8'h00;
    mem['h463C]=8'h00; mem['h463D]=8'h00; mem['h463E]=8'h00; mem['h463F]=8'h00;
    mem['h4640]=8'h00; mem['h4641]=8'h00; mem['h4642]=8'h00; mem['h4643]=8'h00;
    mem['h4644]=8'h00; mem['h4645]=8'h00; mem['h4646]=8'h00; mem['h4647]=8'h00;
    mem['h4648]=8'h00; mem['h4649]=8'h00; mem['h464A]=8'h00; mem['h464B]=8'h00;
    mem['h464C]=8'h00; mem['h464D]=8'h00; mem['h464E]=8'h00; mem['h464F]=8'h00;
    mem['h4650]=8'h00; mem['h4651]=8'h00; mem['h4652]=8'h00; mem['h4653]=8'h00;
    mem['h4654]=8'h00; mem['h4655]=8'h00; mem['h4656]=8'h00; mem['h4657]=8'h00;
    mem['h4658]=8'h00; mem['h4659]=8'h00; mem['h465A]=8'h00; mem['h465B]=8'h00;
    mem['h465C]=8'h00; mem['h465D]=8'h00; mem['h465E]=8'h00; mem['h465F]=8'h00;
    mem['h4660]=8'h00; mem['h4661]=8'h00; mem['h4662]=8'h00; mem['h4663]=8'h00;
    mem['h4664]=8'h00; mem['h4665]=8'h00; mem['h4666]=8'h00; mem['h4667]=8'h00;
    mem['h4668]=8'h00; mem['h4669]=8'h00; mem['h466A]=8'h00; mem['h466B]=8'h00;
    mem['h466C]=8'h00; mem['h466D]=8'h00; mem['h466E]=8'h00; mem['h466F]=8'h00;
    mem['h4670]=8'h00; mem['h4671]=8'h00; mem['h4672]=8'h00; mem['h4673]=8'h00;
    mem['h4674]=8'h00; mem['h4675]=8'h00; mem['h4676]=8'h00; mem['h4677]=8'h00;
    mem['h4678]=8'h00; mem['h4679]=8'h00; mem['h467A]=8'h00; mem['h467B]=8'h00;
    mem['h467C]=8'h00; mem['h467D]=8'h00; mem['h467E]=8'h00; mem['h467F]=8'h00;
    mem['h4680]=8'h00; mem['h4681]=8'h00; mem['h4682]=8'h00; mem['h4683]=8'h00;
    mem['h4684]=8'h00; mem['h4685]=8'h00; mem['h4686]=8'h00; mem['h4687]=8'h00;
    mem['h4688]=8'h00; mem['h4689]=8'h00; mem['h468A]=8'h00; mem['h468B]=8'h00;
    mem['h468C]=8'h00; mem['h468D]=8'h00; mem['h468E]=8'h00; mem['h468F]=8'h00;
    mem['h4690]=8'h00; mem['h4691]=8'h00; mem['h4692]=8'h00; mem['h4693]=8'h00;
    mem['h4694]=8'h00; mem['h4695]=8'h00; mem['h4696]=8'h00; mem['h4697]=8'h00;
    mem['h4698]=8'h00; mem['h4699]=8'h00; mem['h469A]=8'h00; mem['h469B]=8'h00;
    mem['h469C]=8'h00; mem['h469D]=8'h00; mem['h469E]=8'h00; mem['h469F]=8'h00;
    mem['h46A0]=8'h00; mem['h46A1]=8'h00; mem['h46A2]=8'h00; mem['h46A3]=8'h00;
    mem['h46A4]=8'h00; mem['h46A5]=8'h00; mem['h46A6]=8'h00; mem['h46A7]=8'h00;
    mem['h46A8]=8'h00; mem['h46A9]=8'h00; mem['h46AA]=8'h00; mem['h46AB]=8'h00;
    mem['h46AC]=8'h00; mem['h46AD]=8'h00; mem['h46AE]=8'h00; mem['h46AF]=8'h00;
    mem['h46B0]=8'h00; mem['h46B1]=8'h00; mem['h46B2]=8'h00; mem['h46B3]=8'h00;
    mem['h46B4]=8'h00; mem['h46B5]=8'h00; mem['h46B6]=8'h00; mem['h46B7]=8'h00;
    mem['h46B8]=8'h00; mem['h46B9]=8'h00; mem['h46BA]=8'h00; mem['h46BB]=8'h00;
    mem['h46BC]=8'h00; mem['h46BD]=8'h00; mem['h46BE]=8'h00; mem['h46BF]=8'h00;
    mem['h46C0]=8'h00; mem['h46C1]=8'h00; mem['h46C2]=8'h00; mem['h46C3]=8'h00;
    mem['h46C4]=8'h00; mem['h46C5]=8'h00; mem['h46C6]=8'h00; mem['h46C7]=8'h00;
    mem['h46C8]=8'h00; mem['h46C9]=8'h00; mem['h46CA]=8'h00; mem['h46CB]=8'h00;
    mem['h46CC]=8'h00; mem['h46CD]=8'h00; mem['h46CE]=8'h00; mem['h46CF]=8'h00;
    mem['h46D0]=8'h00; mem['h46D1]=8'h00; mem['h46D2]=8'h00; mem['h46D3]=8'h00;
    mem['h46D4]=8'h00; mem['h46D5]=8'h00; mem['h46D6]=8'h00; mem['h46D7]=8'h00;
    mem['h46D8]=8'h00; mem['h46D9]=8'h00; mem['h46DA]=8'h00; mem['h46DB]=8'h00;
    mem['h46DC]=8'h00; mem['h46DD]=8'h00; mem['h46DE]=8'h00; mem['h46DF]=8'h00;
    mem['h46E0]=8'h00; mem['h46E1]=8'h00; mem['h46E2]=8'h00; mem['h46E3]=8'h00;
    mem['h46E4]=8'h00; mem['h46E5]=8'h00; mem['h46E6]=8'h00; mem['h46E7]=8'h00;
    mem['h46E8]=8'h00; mem['h46E9]=8'h00; mem['h46EA]=8'h00; mem['h46EB]=8'h00;
    mem['h46EC]=8'h00; mem['h46ED]=8'h00; mem['h46EE]=8'h00; mem['h46EF]=8'h00;
    mem['h46F0]=8'h00; mem['h46F1]=8'h00; mem['h46F2]=8'h00; mem['h46F3]=8'h00;
    mem['h46F4]=8'h00; mem['h46F5]=8'h00; mem['h46F6]=8'h00; mem['h46F7]=8'h00;
    mem['h46F8]=8'h00; mem['h46F9]=8'h00; mem['h46FA]=8'h00; mem['h46FB]=8'h00;
    mem['h46FC]=8'h00; mem['h46FD]=8'h00; mem['h46FE]=8'h00; mem['h46FF]=8'h00;
    mem['h4700]=8'h00; mem['h4701]=8'h00; mem['h4702]=8'h00; mem['h4703]=8'h00;
    mem['h4704]=8'h00; mem['h4705]=8'h00; mem['h4706]=8'h00; mem['h4707]=8'h00;
    mem['h4708]=8'h00; mem['h4709]=8'h00; mem['h470A]=8'h00; mem['h470B]=8'h00;
    mem['h470C]=8'h00; mem['h470D]=8'h00; mem['h470E]=8'h00; mem['h470F]=8'h00;
    mem['h4710]=8'h00; mem['h4711]=8'h00; mem['h4712]=8'h00; mem['h4713]=8'h00;
    mem['h4714]=8'h00; mem['h4715]=8'h00; mem['h4716]=8'h00; mem['h4717]=8'h00;
    mem['h4718]=8'h00; mem['h4719]=8'h00; mem['h471A]=8'h00; mem['h471B]=8'h00;
    mem['h471C]=8'h00; mem['h471D]=8'h00; mem['h471E]=8'h00; mem['h471F]=8'h00;
    mem['h4720]=8'h00; mem['h4721]=8'h00; mem['h4722]=8'h00; mem['h4723]=8'h00;
    mem['h4724]=8'h00; mem['h4725]=8'h00; mem['h4726]=8'h00; mem['h4727]=8'h00;
    mem['h4728]=8'h00; mem['h4729]=8'h00; mem['h472A]=8'h00; mem['h472B]=8'h00;
    mem['h472C]=8'h00; mem['h472D]=8'h00; mem['h472E]=8'h00; mem['h472F]=8'h00;
    mem['h4730]=8'h00; mem['h4731]=8'h00; mem['h4732]=8'h00; mem['h4733]=8'h00;
    mem['h4734]=8'h00; mem['h4735]=8'h00; mem['h4736]=8'h00; mem['h4737]=8'h00;
    mem['h4738]=8'h00; mem['h4739]=8'h00; mem['h473A]=8'h00; mem['h473B]=8'h00;
    mem['h473C]=8'h00; mem['h473D]=8'h00; mem['h473E]=8'h00; mem['h473F]=8'h00;
    mem['h4740]=8'h00; mem['h4741]=8'h00; mem['h4742]=8'h00; mem['h4743]=8'h00;
    mem['h4744]=8'h00; mem['h4745]=8'h00; mem['h4746]=8'h00; mem['h4747]=8'h00;
    mem['h4748]=8'h00; mem['h4749]=8'h00; mem['h474A]=8'h00; mem['h474B]=8'h00;
    mem['h474C]=8'h00; mem['h474D]=8'h00; mem['h474E]=8'h00; mem['h474F]=8'h00;
    mem['h4750]=8'h00; mem['h4751]=8'h00; mem['h4752]=8'h00; mem['h4753]=8'h00;
    mem['h4754]=8'h00; mem['h4755]=8'h00; mem['h4756]=8'h00; mem['h4757]=8'h00;
    mem['h4758]=8'h00; mem['h4759]=8'h00; mem['h475A]=8'h00; mem['h475B]=8'h00;
    mem['h475C]=8'h00; mem['h475D]=8'h00; mem['h475E]=8'h00; mem['h475F]=8'h00;
    mem['h4760]=8'h00; mem['h4761]=8'h00; mem['h4762]=8'h00; mem['h4763]=8'h00;
    mem['h4764]=8'h00; mem['h4765]=8'h00; mem['h4766]=8'h00; mem['h4767]=8'h00;
    mem['h4768]=8'h00; mem['h4769]=8'h00; mem['h476A]=8'h00; mem['h476B]=8'h00;
    mem['h476C]=8'h00; mem['h476D]=8'h00; mem['h476E]=8'h00; mem['h476F]=8'h00;
    mem['h4770]=8'h00; mem['h4771]=8'h00; mem['h4772]=8'h00; mem['h4773]=8'h00;
    mem['h4774]=8'h00; mem['h4775]=8'h00; mem['h4776]=8'h00; mem['h4777]=8'h00;
    mem['h4778]=8'h00; mem['h4779]=8'h00; mem['h477A]=8'h00; mem['h477B]=8'h00;
    mem['h477C]=8'h00; mem['h477D]=8'h00; mem['h477E]=8'h00; mem['h477F]=8'h00;
    mem['h4780]=8'h00; mem['h4781]=8'h00; mem['h4782]=8'h00; mem['h4783]=8'h00;
    mem['h4784]=8'h00; mem['h4785]=8'h00; mem['h4786]=8'h00; mem['h4787]=8'h00;
    mem['h4788]=8'h00; mem['h4789]=8'h00; mem['h478A]=8'h00; mem['h478B]=8'h00;
    mem['h478C]=8'h00; mem['h478D]=8'h00; mem['h478E]=8'h00; mem['h478F]=8'h00;
    mem['h4790]=8'h00; mem['h4791]=8'h00; mem['h4792]=8'h00; mem['h4793]=8'h00;
    mem['h4794]=8'h00; mem['h4795]=8'h00; mem['h4796]=8'h00; mem['h4797]=8'h00;
    mem['h4798]=8'h00; mem['h4799]=8'h00; mem['h479A]=8'h00; mem['h479B]=8'h00;
    mem['h479C]=8'h00; mem['h479D]=8'h00; mem['h479E]=8'h00; mem['h479F]=8'h00;
    mem['h47A0]=8'h00; mem['h47A1]=8'h00; mem['h47A2]=8'h00; mem['h47A3]=8'h00;
    mem['h47A4]=8'h00; mem['h47A5]=8'h00; mem['h47A6]=8'h00; mem['h47A7]=8'h00;
    mem['h47A8]=8'h00; mem['h47A9]=8'h00; mem['h47AA]=8'h00; mem['h47AB]=8'h00;
    mem['h47AC]=8'h00; mem['h47AD]=8'h00; mem['h47AE]=8'h00; mem['h47AF]=8'h00;
    mem['h47B0]=8'h00; mem['h47B1]=8'h00; mem['h47B2]=8'h00; mem['h47B3]=8'h00;
    mem['h47B4]=8'h00; mem['h47B5]=8'h00; mem['h47B6]=8'h00; mem['h47B7]=8'h00;
    mem['h47B8]=8'h00; mem['h47B9]=8'h00; mem['h47BA]=8'h00; mem['h47BB]=8'h00;
    mem['h47BC]=8'h00; mem['h47BD]=8'h00; mem['h47BE]=8'h00; mem['h47BF]=8'h00;
    mem['h47C0]=8'h00; mem['h47C1]=8'h00; mem['h47C2]=8'h00; mem['h47C3]=8'h00;
    mem['h47C4]=8'h00; mem['h47C5]=8'h00; mem['h47C6]=8'h00; mem['h47C7]=8'h00;
    mem['h47C8]=8'h00; mem['h47C9]=8'h00; mem['h47CA]=8'h00; mem['h47CB]=8'h00;
    mem['h47CC]=8'h00; mem['h47CD]=8'h00; mem['h47CE]=8'h00; mem['h47CF]=8'h00;
    mem['h47D0]=8'h00; mem['h47D1]=8'h00; mem['h47D2]=8'h00; mem['h47D3]=8'h00;
    mem['h47D4]=8'h00; mem['h47D5]=8'h00; mem['h47D6]=8'h00; mem['h47D7]=8'h00;
    mem['h47D8]=8'h00; mem['h47D9]=8'h00; mem['h47DA]=8'h00; mem['h47DB]=8'h00;
    mem['h47DC]=8'h00; mem['h47DD]=8'h00; mem['h47DE]=8'h00; mem['h47DF]=8'h00;
    mem['h47E0]=8'h00; mem['h47E1]=8'h00; mem['h47E2]=8'h00; mem['h47E3]=8'h00;
    mem['h47E4]=8'h00; mem['h47E5]=8'h00; mem['h47E6]=8'h00; mem['h47E7]=8'h00;
    mem['h47E8]=8'h00; mem['h47E9]=8'h00; mem['h47EA]=8'h00; mem['h47EB]=8'h00;
    mem['h47EC]=8'h00; mem['h47ED]=8'h00; mem['h47EE]=8'h00; mem['h47EF]=8'h00;
    mem['h47F0]=8'h00; mem['h47F1]=8'h00; mem['h47F2]=8'h00; mem['h47F3]=8'h00;
    mem['h47F4]=8'h00; mem['h47F5]=8'h00; mem['h47F6]=8'h00; mem['h47F7]=8'h00;
    mem['h47F8]=8'h00; mem['h47F9]=8'h00; mem['h47FA]=8'h00; mem['h47FB]=8'h00;
    mem['h47FC]=8'h00; mem['h47FD]=8'h00; mem['h47FE]=8'h00; mem['h47FF]=8'h00;
    mem['h4800]=8'h00; mem['h4801]=8'h00; mem['h4802]=8'h00; mem['h4803]=8'h00;
    mem['h4804]=8'h00; mem['h4805]=8'h00; mem['h4806]=8'h00; mem['h4807]=8'h00;
    mem['h4808]=8'h00; mem['h4809]=8'h00; mem['h480A]=8'h00; mem['h480B]=8'h00;
    mem['h480C]=8'h00; mem['h480D]=8'h00; mem['h480E]=8'h00; mem['h480F]=8'h00;
    mem['h4810]=8'h00; mem['h4811]=8'h00; mem['h4812]=8'h00; mem['h4813]=8'h00;
    mem['h4814]=8'h00; mem['h4815]=8'h00; mem['h4816]=8'h00; mem['h4817]=8'h00;
    mem['h4818]=8'h00; mem['h4819]=8'h00; mem['h481A]=8'h00; mem['h481B]=8'h00;
    mem['h481C]=8'h00; mem['h481D]=8'h00; mem['h481E]=8'h00; mem['h481F]=8'h00;
    mem['h4820]=8'h00; mem['h4821]=8'h00; mem['h4822]=8'h00; mem['h4823]=8'h00;
    mem['h4824]=8'h00; mem['h4825]=8'h00; mem['h4826]=8'h00; mem['h4827]=8'h00;
    mem['h4828]=8'h00; mem['h4829]=8'h00; mem['h482A]=8'h00; mem['h482B]=8'h00;
    mem['h482C]=8'h00; mem['h482D]=8'h00; mem['h482E]=8'h00; mem['h482F]=8'h00;
    mem['h4830]=8'h00; mem['h4831]=8'h00; mem['h4832]=8'h00; mem['h4833]=8'h00;
    mem['h4834]=8'h00; mem['h4835]=8'h00; mem['h4836]=8'h00; mem['h4837]=8'h00;
    mem['h4838]=8'h00; mem['h4839]=8'h00; mem['h483A]=8'h00; mem['h483B]=8'h00;
    mem['h483C]=8'h00; mem['h483D]=8'h00; mem['h483E]=8'h00; mem['h483F]=8'h00;
    mem['h4840]=8'h00; mem['h4841]=8'h00; mem['h4842]=8'h00; mem['h4843]=8'h00;
    mem['h4844]=8'h00; mem['h4845]=8'h00; mem['h4846]=8'h00; mem['h4847]=8'h00;
    mem['h4848]=8'h00; mem['h4849]=8'h00; mem['h484A]=8'h00; mem['h484B]=8'h00;
    mem['h484C]=8'h00; mem['h484D]=8'h00; mem['h484E]=8'h00; mem['h484F]=8'h00;
    mem['h4850]=8'h00; mem['h4851]=8'h00; mem['h4852]=8'h00; mem['h4853]=8'h00;
    mem['h4854]=8'h00; mem['h4855]=8'h00; mem['h4856]=8'h00; mem['h4857]=8'h00;
    mem['h4858]=8'h00; mem['h4859]=8'h00; mem['h485A]=8'h00; mem['h485B]=8'h00;
    mem['h485C]=8'h00; mem['h485D]=8'h00; mem['h485E]=8'h00; mem['h485F]=8'h00;
    mem['h4860]=8'h00; mem['h4861]=8'h00; mem['h4862]=8'h00; mem['h4863]=8'h00;
    mem['h4864]=8'h00; mem['h4865]=8'h00; mem['h4866]=8'h00; mem['h4867]=8'h00;
    mem['h4868]=8'h00; mem['h4869]=8'h00; mem['h486A]=8'h00; mem['h486B]=8'h00;
    mem['h486C]=8'h00; mem['h486D]=8'h00; mem['h486E]=8'h00; mem['h486F]=8'h00;
    mem['h4870]=8'h00; mem['h4871]=8'h00; mem['h4872]=8'h00; mem['h4873]=8'h00;
    mem['h4874]=8'h00; mem['h4875]=8'h00; mem['h4876]=8'h00; mem['h4877]=8'h00;
    mem['h4878]=8'h00; mem['h4879]=8'h00; mem['h487A]=8'h00; mem['h487B]=8'h00;
    mem['h487C]=8'h00; mem['h487D]=8'h00; mem['h487E]=8'h00; mem['h487F]=8'h00;
    mem['h4880]=8'h00; mem['h4881]=8'h00; mem['h4882]=8'h00; mem['h4883]=8'h00;
    mem['h4884]=8'h00; mem['h4885]=8'h00; mem['h4886]=8'h00; mem['h4887]=8'h00;
    mem['h4888]=8'h00; mem['h4889]=8'h00; mem['h488A]=8'h00; mem['h488B]=8'h00;
    mem['h488C]=8'h00; mem['h488D]=8'h00; mem['h488E]=8'h00; mem['h488F]=8'h00;
    mem['h4890]=8'h00; mem['h4891]=8'h00; mem['h4892]=8'h00; mem['h4893]=8'h00;
    mem['h4894]=8'h00; mem['h4895]=8'h00; mem['h4896]=8'h00; mem['h4897]=8'h00;
    mem['h4898]=8'h00; mem['h4899]=8'h00; mem['h489A]=8'h00; mem['h489B]=8'h00;
    mem['h489C]=8'h00; mem['h489D]=8'h00; mem['h489E]=8'h00; mem['h489F]=8'h00;
    mem['h48A0]=8'h00; mem['h48A1]=8'h00; mem['h48A2]=8'h00; mem['h48A3]=8'h00;
    mem['h48A4]=8'h00; mem['h48A5]=8'h00; mem['h48A6]=8'h00; mem['h48A7]=8'h00;
    mem['h48A8]=8'h00; mem['h48A9]=8'h00; mem['h48AA]=8'h00; mem['h48AB]=8'h00;
    mem['h48AC]=8'h00; mem['h48AD]=8'h00; mem['h48AE]=8'h00; mem['h48AF]=8'h00;
    mem['h48B0]=8'h00; mem['h48B1]=8'h00; mem['h48B2]=8'h00; mem['h48B3]=8'h00;
    mem['h48B4]=8'h00; mem['h48B5]=8'h00; mem['h48B6]=8'h00; mem['h48B7]=8'h00;
    mem['h48B8]=8'h00; mem['h48B9]=8'h00; mem['h48BA]=8'h00; mem['h48BB]=8'h00;
    mem['h48BC]=8'h00; mem['h48BD]=8'h00; mem['h48BE]=8'h00; mem['h48BF]=8'h00;
    mem['h48C0]=8'h00; mem['h48C1]=8'h00; mem['h48C2]=8'h00; mem['h48C3]=8'h00;
    mem['h48C4]=8'h00; mem['h48C5]=8'h00; mem['h48C6]=8'h00; mem['h48C7]=8'h00;
    mem['h48C8]=8'h00; mem['h48C9]=8'h00; mem['h48CA]=8'h00; mem['h48CB]=8'h00;
    mem['h48CC]=8'h00; mem['h48CD]=8'h00; mem['h48CE]=8'h00; mem['h48CF]=8'h00;
    mem['h48D0]=8'h00; mem['h48D1]=8'h00; mem['h48D2]=8'h00; mem['h48D3]=8'h00;
    mem['h48D4]=8'h00; mem['h48D5]=8'h00; mem['h48D6]=8'h00; mem['h48D7]=8'h00;
    mem['h48D8]=8'h00; mem['h48D9]=8'h00; mem['h48DA]=8'h00; mem['h48DB]=8'h00;
    mem['h48DC]=8'h00; mem['h48DD]=8'h00; mem['h48DE]=8'h00; mem['h48DF]=8'h00;
    mem['h48E0]=8'h00; mem['h48E1]=8'h00; mem['h48E2]=8'h00; mem['h48E3]=8'h00;
    mem['h48E4]=8'h00; mem['h48E5]=8'h00; mem['h48E6]=8'h00; mem['h48E7]=8'h00;
    mem['h48E8]=8'h00; mem['h48E9]=8'h00; mem['h48EA]=8'h00; mem['h48EB]=8'h00;
    mem['h48EC]=8'h00; mem['h48ED]=8'h00; mem['h48EE]=8'h00; mem['h48EF]=8'h00;
    mem['h48F0]=8'h00; mem['h48F1]=8'h00; mem['h48F2]=8'h00; mem['h48F3]=8'h00;
    mem['h48F4]=8'h00; mem['h48F5]=8'h00; mem['h48F6]=8'h00; mem['h48F7]=8'h00;
    mem['h48F8]=8'h00; mem['h48F9]=8'h00; mem['h48FA]=8'h00; mem['h48FB]=8'h00;
    mem['h48FC]=8'h00; mem['h48FD]=8'h00; mem['h48FE]=8'h00; mem['h48FF]=8'h00;
    mem['h4900]=8'h00; mem['h4901]=8'h00; mem['h4902]=8'h00; mem['h4903]=8'h00;
    mem['h4904]=8'h00; mem['h4905]=8'h00; mem['h4906]=8'h00; mem['h4907]=8'h00;
    mem['h4908]=8'h00; mem['h4909]=8'h00; mem['h490A]=8'h00; mem['h490B]=8'h00;
    mem['h490C]=8'h00; mem['h490D]=8'h00; mem['h490E]=8'h00; mem['h490F]=8'h00;
    mem['h4910]=8'h00; mem['h4911]=8'h00; mem['h4912]=8'h00; mem['h4913]=8'h00;
    mem['h4914]=8'h00; mem['h4915]=8'h00; mem['h4916]=8'h00; mem['h4917]=8'h00;
    mem['h4918]=8'h00; mem['h4919]=8'h00; mem['h491A]=8'h00; mem['h491B]=8'h00;
    mem['h491C]=8'h00; mem['h491D]=8'h00; mem['h491E]=8'h00; mem['h491F]=8'h00;
    mem['h4920]=8'h00; mem['h4921]=8'h00; mem['h4922]=8'h00; mem['h4923]=8'h00;
    mem['h4924]=8'h00; mem['h4925]=8'h00; mem['h4926]=8'h00; mem['h4927]=8'h00;
    mem['h4928]=8'h00; mem['h4929]=8'h00; mem['h492A]=8'h00; mem['h492B]=8'h00;
    mem['h492C]=8'h00; mem['h492D]=8'h00; mem['h492E]=8'h00; mem['h492F]=8'h00;
    mem['h4930]=8'h00; mem['h4931]=8'h00; mem['h4932]=8'h00; mem['h4933]=8'h00;
    mem['h4934]=8'h00; mem['h4935]=8'h00; mem['h4936]=8'h00; mem['h4937]=8'h00;
    mem['h4938]=8'h00; mem['h4939]=8'h00; mem['h493A]=8'h00; mem['h493B]=8'h00;
    mem['h493C]=8'h00; mem['h493D]=8'h00; mem['h493E]=8'h00; mem['h493F]=8'h00;
    mem['h4940]=8'h00; mem['h4941]=8'h00; mem['h4942]=8'h00; mem['h4943]=8'h00;
    mem['h4944]=8'h00; mem['h4945]=8'h00; mem['h4946]=8'h00; mem['h4947]=8'h00;
    mem['h4948]=8'h00; mem['h4949]=8'h00; mem['h494A]=8'h00; mem['h494B]=8'h00;
    mem['h494C]=8'h00; mem['h494D]=8'h00; mem['h494E]=8'h00; mem['h494F]=8'h00;
    mem['h4950]=8'h00; mem['h4951]=8'h00; mem['h4952]=8'h00; mem['h4953]=8'h00;
    mem['h4954]=8'h00; mem['h4955]=8'h00; mem['h4956]=8'h00; mem['h4957]=8'h00;
    mem['h4958]=8'h00; mem['h4959]=8'h00; mem['h495A]=8'h00; mem['h495B]=8'h00;
    mem['h495C]=8'h00; mem['h495D]=8'h00; mem['h495E]=8'h00; mem['h495F]=8'h00;
    mem['h4960]=8'h00; mem['h4961]=8'h00; mem['h4962]=8'h00; mem['h4963]=8'h00;
    mem['h4964]=8'h00; mem['h4965]=8'h00; mem['h4966]=8'h00; mem['h4967]=8'h00;
    mem['h4968]=8'h00; mem['h4969]=8'h00; mem['h496A]=8'h00; mem['h496B]=8'h00;
    mem['h496C]=8'h00; mem['h496D]=8'h00; mem['h496E]=8'h00; mem['h496F]=8'h00;
    mem['h4970]=8'h00; mem['h4971]=8'h00; mem['h4972]=8'h00; mem['h4973]=8'h00;
    mem['h4974]=8'h00; mem['h4975]=8'h00; mem['h4976]=8'h00; mem['h4977]=8'h00;
    mem['h4978]=8'h00; mem['h4979]=8'h00; mem['h497A]=8'h00; mem['h497B]=8'h00;
    mem['h497C]=8'h00; mem['h497D]=8'h00; mem['h497E]=8'h00; mem['h497F]=8'h00;
    mem['h4980]=8'h00; mem['h4981]=8'h00; mem['h4982]=8'h00; mem['h4983]=8'h00;
    mem['h4984]=8'h00; mem['h4985]=8'h00; mem['h4986]=8'h00; mem['h4987]=8'h00;
    mem['h4988]=8'h00; mem['h4989]=8'h00; mem['h498A]=8'h00; mem['h498B]=8'h00;
    mem['h498C]=8'h00; mem['h498D]=8'h00; mem['h498E]=8'h00; mem['h498F]=8'h00;
    mem['h4990]=8'h00; mem['h4991]=8'h00; mem['h4992]=8'h00; mem['h4993]=8'h00;
    mem['h4994]=8'h00; mem['h4995]=8'h00; mem['h4996]=8'h00; mem['h4997]=8'h00;
    mem['h4998]=8'h00; mem['h4999]=8'h00; mem['h499A]=8'h00; mem['h499B]=8'h00;
    mem['h499C]=8'h00; mem['h499D]=8'h00; mem['h499E]=8'h00; mem['h499F]=8'h00;
    mem['h49A0]=8'h00; mem['h49A1]=8'h00; mem['h49A2]=8'h00; mem['h49A3]=8'h00;
    mem['h49A4]=8'h00; mem['h49A5]=8'h00; mem['h49A6]=8'h00; mem['h49A7]=8'h00;
    mem['h49A8]=8'h00; mem['h49A9]=8'h00; mem['h49AA]=8'h00; mem['h49AB]=8'h00;
    mem['h49AC]=8'h00; mem['h49AD]=8'h00; mem['h49AE]=8'h00; mem['h49AF]=8'h00;
    mem['h49B0]=8'h00; mem['h49B1]=8'h00; mem['h49B2]=8'h00; mem['h49B3]=8'h00;
    mem['h49B4]=8'h00; mem['h49B5]=8'h00; mem['h49B6]=8'h00; mem['h49B7]=8'h00;
    mem['h49B8]=8'h00; mem['h49B9]=8'h00; mem['h49BA]=8'h00; mem['h49BB]=8'h00;
    mem['h49BC]=8'h00; mem['h49BD]=8'h00; mem['h49BE]=8'h00; mem['h49BF]=8'h00;
    mem['h49C0]=8'h00; mem['h49C1]=8'h00; mem['h49C2]=8'h00; mem['h49C3]=8'h00;
    mem['h49C4]=8'h00; mem['h49C5]=8'h00; mem['h49C6]=8'h00; mem['h49C7]=8'h00;
    mem['h49C8]=8'h00; mem['h49C9]=8'h00; mem['h49CA]=8'h00; mem['h49CB]=8'h00;
    mem['h49CC]=8'h00; mem['h49CD]=8'h00; mem['h49CE]=8'h00; mem['h49CF]=8'h00;
    mem['h49D0]=8'h00; mem['h49D1]=8'h00; mem['h49D2]=8'h00; mem['h49D3]=8'h00;
    mem['h49D4]=8'h00; mem['h49D5]=8'h00; mem['h49D6]=8'h00; mem['h49D7]=8'h00;
    mem['h49D8]=8'h00; mem['h49D9]=8'h00; mem['h49DA]=8'h00; mem['h49DB]=8'h00;
    mem['h49DC]=8'h00; mem['h49DD]=8'h00; mem['h49DE]=8'h00; mem['h49DF]=8'h00;
    mem['h49E0]=8'h00; mem['h49E1]=8'h00; mem['h49E2]=8'h00; mem['h49E3]=8'h00;
    mem['h49E4]=8'h00; mem['h49E5]=8'h00; mem['h49E6]=8'h00; mem['h49E7]=8'h00;
    mem['h49E8]=8'h00; mem['h49E9]=8'h00; mem['h49EA]=8'h00; mem['h49EB]=8'h00;
    mem['h49EC]=8'h00; mem['h49ED]=8'h00; mem['h49EE]=8'h00; mem['h49EF]=8'h00;
    mem['h49F0]=8'h00; mem['h49F1]=8'h00; mem['h49F2]=8'h00; mem['h49F3]=8'h00;
    mem['h49F4]=8'h00; mem['h49F5]=8'h00; mem['h49F6]=8'h00; mem['h49F7]=8'h00;
    mem['h49F8]=8'h00; mem['h49F9]=8'h00; mem['h49FA]=8'h00; mem['h49FB]=8'h00;
    mem['h49FC]=8'h00; mem['h49FD]=8'h00; mem['h49FE]=8'h00; mem['h49FF]=8'h00;
    mem['h4A00]=8'h00; mem['h4A01]=8'h00; mem['h4A02]=8'h00; mem['h4A03]=8'h00;
    mem['h4A04]=8'h00; mem['h4A05]=8'h00; mem['h4A06]=8'h00; mem['h4A07]=8'h00;
    mem['h4A08]=8'h00; mem['h4A09]=8'h00; mem['h4A0A]=8'h00; mem['h4A0B]=8'h00;
    mem['h4A0C]=8'h00; mem['h4A0D]=8'h00; mem['h4A0E]=8'h00; mem['h4A0F]=8'h00;
    mem['h4A10]=8'h00; mem['h4A11]=8'h00; mem['h4A12]=8'h00; mem['h4A13]=8'h00;
    mem['h4A14]=8'h00; mem['h4A15]=8'h00; mem['h4A16]=8'h00; mem['h4A17]=8'h00;
    mem['h4A18]=8'h00; mem['h4A19]=8'h00; mem['h4A1A]=8'h00; mem['h4A1B]=8'h00;
    mem['h4A1C]=8'h00; mem['h4A1D]=8'h00; mem['h4A1E]=8'h00; mem['h4A1F]=8'h00;
    mem['h4A20]=8'h00; mem['h4A21]=8'h00; mem['h4A22]=8'h00; mem['h4A23]=8'h00;
    mem['h4A24]=8'h00; mem['h4A25]=8'h00; mem['h4A26]=8'h00; mem['h4A27]=8'h00;
    mem['h4A28]=8'h00; mem['h4A29]=8'h00; mem['h4A2A]=8'h00; mem['h4A2B]=8'h00;
    mem['h4A2C]=8'h00; mem['h4A2D]=8'h00; mem['h4A2E]=8'h00; mem['h4A2F]=8'h00;
    mem['h4A30]=8'h00; mem['h4A31]=8'h00; mem['h4A32]=8'h00; mem['h4A33]=8'h00;
    mem['h4A34]=8'h00; mem['h4A35]=8'h00; mem['h4A36]=8'h00; mem['h4A37]=8'h00;
    mem['h4A38]=8'h00; mem['h4A39]=8'h00; mem['h4A3A]=8'h00; mem['h4A3B]=8'h00;
    mem['h4A3C]=8'h00; mem['h4A3D]=8'h00; mem['h4A3E]=8'h00; mem['h4A3F]=8'h00;
    mem['h4A40]=8'h00; mem['h4A41]=8'h00; mem['h4A42]=8'h00; mem['h4A43]=8'h00;
    mem['h4A44]=8'h00; mem['h4A45]=8'h00; mem['h4A46]=8'h00; mem['h4A47]=8'h00;
    mem['h4A48]=8'h00; mem['h4A49]=8'h00; mem['h4A4A]=8'h00; mem['h4A4B]=8'h00;
    mem['h4A4C]=8'h00; mem['h4A4D]=8'h00; mem['h4A4E]=8'h00; mem['h4A4F]=8'h00;
    mem['h4A50]=8'h00; mem['h4A51]=8'h00; mem['h4A52]=8'h00; mem['h4A53]=8'h00;
    mem['h4A54]=8'h00; mem['h4A55]=8'h00; mem['h4A56]=8'h00; mem['h4A57]=8'h00;
    mem['h4A58]=8'h00; mem['h4A59]=8'h00; mem['h4A5A]=8'h00; mem['h4A5B]=8'h00;
    mem['h4A5C]=8'h00; mem['h4A5D]=8'h00; mem['h4A5E]=8'h00; mem['h4A5F]=8'h00;
    mem['h4A60]=8'h00; mem['h4A61]=8'h00; mem['h4A62]=8'h00; mem['h4A63]=8'h00;
    mem['h4A64]=8'h00; mem['h4A65]=8'h00; mem['h4A66]=8'h00; mem['h4A67]=8'h00;
    mem['h4A68]=8'h00; mem['h4A69]=8'h00; mem['h4A6A]=8'h00; mem['h4A6B]=8'h00;
    mem['h4A6C]=8'h00; mem['h4A6D]=8'h00; mem['h4A6E]=8'h00; mem['h4A6F]=8'h00;
    mem['h4A70]=8'h00; mem['h4A71]=8'h00; mem['h4A72]=8'h00; mem['h4A73]=8'h00;
    mem['h4A74]=8'h00; mem['h4A75]=8'h00; mem['h4A76]=8'h00; mem['h4A77]=8'h00;
    mem['h4A78]=8'h00; mem['h4A79]=8'h00; mem['h4A7A]=8'h00; mem['h4A7B]=8'h00;
    mem['h4A7C]=8'h00; mem['h4A7D]=8'h00; mem['h4A7E]=8'h00; mem['h4A7F]=8'h00;
    mem['h4A80]=8'h00; mem['h4A81]=8'h00; mem['h4A82]=8'h00; mem['h4A83]=8'h00;
    mem['h4A84]=8'h00; mem['h4A85]=8'h00; mem['h4A86]=8'h00; mem['h4A87]=8'h00;
    mem['h4A88]=8'h00; mem['h4A89]=8'h00; mem['h4A8A]=8'h00; mem['h4A8B]=8'h00;
    mem['h4A8C]=8'h00; mem['h4A8D]=8'h00; mem['h4A8E]=8'h00; mem['h4A8F]=8'h00;
    mem['h4A90]=8'h00; mem['h4A91]=8'h00; mem['h4A92]=8'h00; mem['h4A93]=8'h00;
    mem['h4A94]=8'h00; mem['h4A95]=8'h00; mem['h4A96]=8'h00; mem['h4A97]=8'h00;
    mem['h4A98]=8'h00; mem['h4A99]=8'h00; mem['h4A9A]=8'h00; mem['h4A9B]=8'h00;
    mem['h4A9C]=8'h00; mem['h4A9D]=8'h00; mem['h4A9E]=8'h00; mem['h4A9F]=8'h00;
    mem['h4AA0]=8'h00; mem['h4AA1]=8'h00; mem['h4AA2]=8'h00; mem['h4AA3]=8'h00;
    mem['h4AA4]=8'h00; mem['h4AA5]=8'h00; mem['h4AA6]=8'h00; mem['h4AA7]=8'h00;
    mem['h4AA8]=8'h00; mem['h4AA9]=8'h00; mem['h4AAA]=8'h00; mem['h4AAB]=8'h00;
    mem['h4AAC]=8'h00; mem['h4AAD]=8'h00; mem['h4AAE]=8'h00; mem['h4AAF]=8'h00;
    mem['h4AB0]=8'h00; mem['h4AB1]=8'h00; mem['h4AB2]=8'h00; mem['h4AB3]=8'h00;
    mem['h4AB4]=8'h00; mem['h4AB5]=8'h00; mem['h4AB6]=8'h00; mem['h4AB7]=8'h00;
    mem['h4AB8]=8'h00; mem['h4AB9]=8'h00; mem['h4ABA]=8'h00; mem['h4ABB]=8'h00;
    mem['h4ABC]=8'h00; mem['h4ABD]=8'h00; mem['h4ABE]=8'h00; mem['h4ABF]=8'h00;
    mem['h4AC0]=8'h00; mem['h4AC1]=8'h00; mem['h4AC2]=8'h00; mem['h4AC3]=8'h00;
    mem['h4AC4]=8'h00; mem['h4AC5]=8'h00; mem['h4AC6]=8'h00; mem['h4AC7]=8'h00;
    mem['h4AC8]=8'h00; mem['h4AC9]=8'h00; mem['h4ACA]=8'h00; mem['h4ACB]=8'h00;
    mem['h4ACC]=8'h00; mem['h4ACD]=8'h00; mem['h4ACE]=8'h00; mem['h4ACF]=8'h00;
    mem['h4AD0]=8'h00; mem['h4AD1]=8'h00; mem['h4AD2]=8'h00; mem['h4AD3]=8'h00;
    mem['h4AD4]=8'h00; mem['h4AD5]=8'h00; mem['h4AD6]=8'h00; mem['h4AD7]=8'h00;
    mem['h4AD8]=8'h00; mem['h4AD9]=8'h00; mem['h4ADA]=8'h00; mem['h4ADB]=8'h00;
    mem['h4ADC]=8'h00; mem['h4ADD]=8'h00; mem['h4ADE]=8'h00; mem['h4ADF]=8'h00;
    mem['h4AE0]=8'h00; mem['h4AE1]=8'h00; mem['h4AE2]=8'h00; mem['h4AE3]=8'h00;
    mem['h4AE4]=8'h00; mem['h4AE5]=8'h00; mem['h4AE6]=8'h00; mem['h4AE7]=8'h00;
    mem['h4AE8]=8'h00; mem['h4AE9]=8'h00; mem['h4AEA]=8'h00; mem['h4AEB]=8'h00;
    mem['h4AEC]=8'h00; mem['h4AED]=8'h00; mem['h4AEE]=8'h00; mem['h4AEF]=8'h00;
    mem['h4AF0]=8'h00; mem['h4AF1]=8'h00; mem['h4AF2]=8'h00; mem['h4AF3]=8'h00;
    mem['h4AF4]=8'h00; mem['h4AF5]=8'h00; mem['h4AF6]=8'h00; mem['h4AF7]=8'h00;
    mem['h4AF8]=8'h00; mem['h4AF9]=8'h00; mem['h4AFA]=8'h00; mem['h4AFB]=8'h00;
    mem['h4AFC]=8'h00; mem['h4AFD]=8'h00; mem['h4AFE]=8'h00; mem['h4AFF]=8'h00;
    mem['h4B00]=8'h00; mem['h4B01]=8'h00; mem['h4B02]=8'h00; mem['h4B03]=8'h00;
    mem['h4B04]=8'h00; mem['h4B05]=8'h00; mem['h4B06]=8'h00; mem['h4B07]=8'h00;
    mem['h4B08]=8'h00; mem['h4B09]=8'h00; mem['h4B0A]=8'h00; mem['h4B0B]=8'h00;
    mem['h4B0C]=8'h00; mem['h4B0D]=8'h00; mem['h4B0E]=8'h00; mem['h4B0F]=8'h00;
    mem['h4B10]=8'h00; mem['h4B11]=8'h00; mem['h4B12]=8'h00; mem['h4B13]=8'h00;
    mem['h4B14]=8'h00; mem['h4B15]=8'h00; mem['h4B16]=8'h00; mem['h4B17]=8'h00;
    mem['h4B18]=8'h00; mem['h4B19]=8'h00; mem['h4B1A]=8'h00; mem['h4B1B]=8'h00;
    mem['h4B1C]=8'h00; mem['h4B1D]=8'h00; mem['h4B1E]=8'h00; mem['h4B1F]=8'h00;
    mem['h4B20]=8'h00; mem['h4B21]=8'h00; mem['h4B22]=8'h00; mem['h4B23]=8'h00;
    mem['h4B24]=8'h00; mem['h4B25]=8'h00; mem['h4B26]=8'h00; mem['h4B27]=8'h00;
    mem['h4B28]=8'h00; mem['h4B29]=8'h00; mem['h4B2A]=8'h00; mem['h4B2B]=8'h00;
    mem['h4B2C]=8'h00; mem['h4B2D]=8'h00; mem['h4B2E]=8'h00; mem['h4B2F]=8'h00;
    mem['h4B30]=8'h00; mem['h4B31]=8'h00; mem['h4B32]=8'h00; mem['h4B33]=8'h00;
    mem['h4B34]=8'h00; mem['h4B35]=8'h00; mem['h4B36]=8'h00; mem['h4B37]=8'h00;
    mem['h4B38]=8'h00; mem['h4B39]=8'h00; mem['h4B3A]=8'h00; mem['h4B3B]=8'h00;
    mem['h4B3C]=8'h00; mem['h4B3D]=8'h00; mem['h4B3E]=8'h00; mem['h4B3F]=8'h00;
    mem['h4B40]=8'h00; mem['h4B41]=8'h00; mem['h4B42]=8'h00; mem['h4B43]=8'h00;
    mem['h4B44]=8'h00; mem['h4B45]=8'h00; mem['h4B46]=8'h00; mem['h4B47]=8'h00;
    mem['h4B48]=8'h00; mem['h4B49]=8'h00; mem['h4B4A]=8'h00; mem['h4B4B]=8'h00;
    mem['h4B4C]=8'h00; mem['h4B4D]=8'h00; mem['h4B4E]=8'h00; mem['h4B4F]=8'h00;
    mem['h4B50]=8'h00; mem['h4B51]=8'h00; mem['h4B52]=8'h00; mem['h4B53]=8'h00;
    mem['h4B54]=8'h00; mem['h4B55]=8'h00; mem['h4B56]=8'h00; mem['h4B57]=8'h00;
    mem['h4B58]=8'h00; mem['h4B59]=8'h00; mem['h4B5A]=8'h00; mem['h4B5B]=8'h00;
    mem['h4B5C]=8'h00; mem['h4B5D]=8'h00; mem['h4B5E]=8'h00; mem['h4B5F]=8'h00;
    mem['h4B60]=8'h00; mem['h4B61]=8'h00; mem['h4B62]=8'h00; mem['h4B63]=8'h00;
    mem['h4B64]=8'h00; mem['h4B65]=8'h00; mem['h4B66]=8'h00; mem['h4B67]=8'h00;
    mem['h4B68]=8'h00; mem['h4B69]=8'h00; mem['h4B6A]=8'h00; mem['h4B6B]=8'h00;
    mem['h4B6C]=8'h00; mem['h4B6D]=8'h00; mem['h4B6E]=8'h00; mem['h4B6F]=8'h00;
    mem['h4B70]=8'h00; mem['h4B71]=8'h00; mem['h4B72]=8'h00; mem['h4B73]=8'h00;
    mem['h4B74]=8'h00; mem['h4B75]=8'h00; mem['h4B76]=8'h00; mem['h4B77]=8'h00;
    mem['h4B78]=8'h00; mem['h4B79]=8'h00; mem['h4B7A]=8'h00; mem['h4B7B]=8'h00;
    mem['h4B7C]=8'h00; mem['h4B7D]=8'h00; mem['h4B7E]=8'h00; mem['h4B7F]=8'h00;
    mem['h4B80]=8'h00; mem['h4B81]=8'h00; mem['h4B82]=8'h00; mem['h4B83]=8'h00;
    mem['h4B84]=8'h00; mem['h4B85]=8'h00; mem['h4B86]=8'h00; mem['h4B87]=8'h00;
    mem['h4B88]=8'h00; mem['h4B89]=8'h00; mem['h4B8A]=8'h00; mem['h4B8B]=8'h00;
    mem['h4B8C]=8'h00; mem['h4B8D]=8'h00; mem['h4B8E]=8'h00; mem['h4B8F]=8'h00;
    mem['h4B90]=8'h00; mem['h4B91]=8'h00; mem['h4B92]=8'h00; mem['h4B93]=8'h00;
    mem['h4B94]=8'h00; mem['h4B95]=8'h00; mem['h4B96]=8'h00; mem['h4B97]=8'h00;
    mem['h4B98]=8'h00; mem['h4B99]=8'h00; mem['h4B9A]=8'h00; mem['h4B9B]=8'h00;
    mem['h4B9C]=8'h00; mem['h4B9D]=8'h00; mem['h4B9E]=8'h00; mem['h4B9F]=8'h00;
    mem['h4BA0]=8'h00; mem['h4BA1]=8'h00; mem['h4BA2]=8'h00; mem['h4BA3]=8'h00;
    mem['h4BA4]=8'h00; mem['h4BA5]=8'h00; mem['h4BA6]=8'h00; mem['h4BA7]=8'h00;
    mem['h4BA8]=8'h00; mem['h4BA9]=8'h00; mem['h4BAA]=8'h00; mem['h4BAB]=8'h00;
    mem['h4BAC]=8'h00; mem['h4BAD]=8'h00; mem['h4BAE]=8'h00; mem['h4BAF]=8'h00;
    mem['h4BB0]=8'h00; mem['h4BB1]=8'h00; mem['h4BB2]=8'h00; mem['h4BB3]=8'h00;
    mem['h4BB4]=8'h00; mem['h4BB5]=8'h00; mem['h4BB6]=8'h00; mem['h4BB7]=8'h00;
    mem['h4BB8]=8'h00; mem['h4BB9]=8'h00; mem['h4BBA]=8'h00; mem['h4BBB]=8'h00;
    mem['h4BBC]=8'h00; mem['h4BBD]=8'h00; mem['h4BBE]=8'h00; mem['h4BBF]=8'h00;
    mem['h4BC0]=8'h00; mem['h4BC1]=8'h00; mem['h4BC2]=8'h00; mem['h4BC3]=8'h00;
    mem['h4BC4]=8'h00; mem['h4BC5]=8'h00; mem['h4BC6]=8'h00; mem['h4BC7]=8'h00;
    mem['h4BC8]=8'h00; mem['h4BC9]=8'h00; mem['h4BCA]=8'h00; mem['h4BCB]=8'h00;
    mem['h4BCC]=8'h00; mem['h4BCD]=8'h00; mem['h4BCE]=8'h00; mem['h4BCF]=8'h00;
    mem['h4BD0]=8'h00; mem['h4BD1]=8'h00; mem['h4BD2]=8'h00; mem['h4BD3]=8'h00;
    mem['h4BD4]=8'h00; mem['h4BD5]=8'h00; mem['h4BD6]=8'h00; mem['h4BD7]=8'h00;
    mem['h4BD8]=8'h00; mem['h4BD9]=8'h00; mem['h4BDA]=8'h00; mem['h4BDB]=8'h00;
    mem['h4BDC]=8'h00; mem['h4BDD]=8'h00; mem['h4BDE]=8'h00; mem['h4BDF]=8'h00;
    mem['h4BE0]=8'h00; mem['h4BE1]=8'h00; mem['h4BE2]=8'h00; mem['h4BE3]=8'h00;
    mem['h4BE4]=8'h00; mem['h4BE5]=8'h00; mem['h4BE6]=8'h00; mem['h4BE7]=8'h00;
    mem['h4BE8]=8'h00; mem['h4BE9]=8'h00; mem['h4BEA]=8'h00; mem['h4BEB]=8'h00;
    mem['h4BEC]=8'h00; mem['h4BED]=8'h00; mem['h4BEE]=8'h00; mem['h4BEF]=8'h00;
    mem['h4BF0]=8'h00; mem['h4BF1]=8'h00; mem['h4BF2]=8'h00; mem['h4BF3]=8'h00;
    mem['h4BF4]=8'h00; mem['h4BF5]=8'h00; mem['h4BF6]=8'h00; mem['h4BF7]=8'h00;
    mem['h4BF8]=8'h00; mem['h4BF9]=8'h00; mem['h4BFA]=8'h00; mem['h4BFB]=8'h00;
    mem['h4BFC]=8'h00; mem['h4BFD]=8'h00; mem['h4BFE]=8'h00; mem['h4BFF]=8'h00;
    mem['h4C00]=8'h00; mem['h4C01]=8'h00; mem['h4C02]=8'h00; mem['h4C03]=8'h00;
    mem['h4C04]=8'h00; mem['h4C05]=8'h00; mem['h4C06]=8'h00; mem['h4C07]=8'h00;
    mem['h4C08]=8'h00; mem['h4C09]=8'h00; mem['h4C0A]=8'h00; mem['h4C0B]=8'h00;
    mem['h4C0C]=8'h00; mem['h4C0D]=8'h00; mem['h4C0E]=8'h00; mem['h4C0F]=8'h00;
    mem['h4C10]=8'h00; mem['h4C11]=8'h00; mem['h4C12]=8'h00; mem['h4C13]=8'h00;
    mem['h4C14]=8'h00; mem['h4C15]=8'h00; mem['h4C16]=8'h00; mem['h4C17]=8'h00;
    mem['h4C18]=8'h00; mem['h4C19]=8'h00; mem['h4C1A]=8'h00; mem['h4C1B]=8'h00;
    mem['h4C1C]=8'h00; mem['h4C1D]=8'h00; mem['h4C1E]=8'h00; mem['h4C1F]=8'h00;
    mem['h4C20]=8'h00; mem['h4C21]=8'h00; mem['h4C22]=8'h00; mem['h4C23]=8'h00;
    mem['h4C24]=8'h00; mem['h4C25]=8'h00; mem['h4C26]=8'h00; mem['h4C27]=8'h00;
    mem['h4C28]=8'h00; mem['h4C29]=8'h00; mem['h4C2A]=8'h00; mem['h4C2B]=8'h00;
    mem['h4C2C]=8'h00; mem['h4C2D]=8'h00; mem['h4C2E]=8'h00; mem['h4C2F]=8'h00;
    mem['h4C30]=8'h00; mem['h4C31]=8'h00; mem['h4C32]=8'h00; mem['h4C33]=8'h00;
    mem['h4C34]=8'h00; mem['h4C35]=8'h00; mem['h4C36]=8'h00; mem['h4C37]=8'h00;
    mem['h4C38]=8'h00; mem['h4C39]=8'h00; mem['h4C3A]=8'h00; mem['h4C3B]=8'h00;
    mem['h4C3C]=8'h00; mem['h4C3D]=8'h00; mem['h4C3E]=8'h00; mem['h4C3F]=8'h00;
    mem['h4C40]=8'h00; mem['h4C41]=8'h00; mem['h4C42]=8'h00; mem['h4C43]=8'h00;
    mem['h4C44]=8'h00; mem['h4C45]=8'h00; mem['h4C46]=8'h00; mem['h4C47]=8'h00;
    mem['h4C48]=8'h00; mem['h4C49]=8'h00; mem['h4C4A]=8'h00; mem['h4C4B]=8'h00;
    mem['h4C4C]=8'h00; mem['h4C4D]=8'h00; mem['h4C4E]=8'h00; mem['h4C4F]=8'h00;
    mem['h4C50]=8'h00; mem['h4C51]=8'h00; mem['h4C52]=8'h00; mem['h4C53]=8'h00;
    mem['h4C54]=8'h00; mem['h4C55]=8'h00; mem['h4C56]=8'h00; mem['h4C57]=8'h00;
    mem['h4C58]=8'h00; mem['h4C59]=8'h00; mem['h4C5A]=8'h00; mem['h4C5B]=8'h00;
    mem['h4C5C]=8'h00; mem['h4C5D]=8'h00; mem['h4C5E]=8'h00; mem['h4C5F]=8'h00;
    mem['h4C60]=8'h00; mem['h4C61]=8'h00; mem['h4C62]=8'h00; mem['h4C63]=8'h00;
    mem['h4C64]=8'h00; mem['h4C65]=8'h00; mem['h4C66]=8'h00; mem['h4C67]=8'h00;
    mem['h4C68]=8'h00; mem['h4C69]=8'h00; mem['h4C6A]=8'h00; mem['h4C6B]=8'h00;
    mem['h4C6C]=8'h00; mem['h4C6D]=8'h00; mem['h4C6E]=8'h00; mem['h4C6F]=8'h00;
    mem['h4C70]=8'h00; mem['h4C71]=8'h00; mem['h4C72]=8'h00; mem['h4C73]=8'h00;
    mem['h4C74]=8'h00; mem['h4C75]=8'h00; mem['h4C76]=8'h00; mem['h4C77]=8'h00;
    mem['h4C78]=8'h00; mem['h4C79]=8'h00; mem['h4C7A]=8'h00; mem['h4C7B]=8'h00;
    mem['h4C7C]=8'h00; mem['h4C7D]=8'h00; mem['h4C7E]=8'h00; mem['h4C7F]=8'h00;
    mem['h4C80]=8'h00; mem['h4C81]=8'h00; mem['h4C82]=8'h00; mem['h4C83]=8'h00;
    mem['h4C84]=8'h00; mem['h4C85]=8'h00; mem['h4C86]=8'h00; mem['h4C87]=8'h00;
    mem['h4C88]=8'h00; mem['h4C89]=8'h00; mem['h4C8A]=8'h00; mem['h4C8B]=8'h00;
    mem['h4C8C]=8'h00; mem['h4C8D]=8'h00; mem['h4C8E]=8'h00; mem['h4C8F]=8'h00;
    mem['h4C90]=8'h00; mem['h4C91]=8'h00; mem['h4C92]=8'h00; mem['h4C93]=8'h00;
    mem['h4C94]=8'h00; mem['h4C95]=8'h00; mem['h4C96]=8'h00; mem['h4C97]=8'h00;
    mem['h4C98]=8'h00; mem['h4C99]=8'h00; mem['h4C9A]=8'h00; mem['h4C9B]=8'h00;
    mem['h4C9C]=8'h00; mem['h4C9D]=8'h00; mem['h4C9E]=8'h00; mem['h4C9F]=8'h00;
    mem['h4CA0]=8'h00; mem['h4CA1]=8'h00; mem['h4CA2]=8'h00; mem['h4CA3]=8'h00;
    mem['h4CA4]=8'h00; mem['h4CA5]=8'h00; mem['h4CA6]=8'h00; mem['h4CA7]=8'h00;
    mem['h4CA8]=8'h00; mem['h4CA9]=8'h00; mem['h4CAA]=8'h00; mem['h4CAB]=8'h00;
    mem['h4CAC]=8'h00; mem['h4CAD]=8'h00; mem['h4CAE]=8'h00; mem['h4CAF]=8'h00;
    mem['h4CB0]=8'h00; mem['h4CB1]=8'h00; mem['h4CB2]=8'h00; mem['h4CB3]=8'h00;
    mem['h4CB4]=8'h00; mem['h4CB5]=8'h00; mem['h4CB6]=8'h00; mem['h4CB7]=8'h00;
    mem['h4CB8]=8'h00; mem['h4CB9]=8'h00; mem['h4CBA]=8'h00; mem['h4CBB]=8'h00;
    mem['h4CBC]=8'h00; mem['h4CBD]=8'h00; mem['h4CBE]=8'h00; mem['h4CBF]=8'h00;
    mem['h4CC0]=8'h00; mem['h4CC1]=8'h00; mem['h4CC2]=8'h00; mem['h4CC3]=8'h00;
    mem['h4CC4]=8'h00; mem['h4CC5]=8'h00; mem['h4CC6]=8'h00; mem['h4CC7]=8'h00;
    mem['h4CC8]=8'h00; mem['h4CC9]=8'h00; mem['h4CCA]=8'h00; mem['h4CCB]=8'h00;
    mem['h4CCC]=8'h00; mem['h4CCD]=8'h00; mem['h4CCE]=8'h00; mem['h4CCF]=8'h00;
    mem['h4CD0]=8'h00; mem['h4CD1]=8'h00; mem['h4CD2]=8'h00; mem['h4CD3]=8'h00;
    mem['h4CD4]=8'h00; mem['h4CD5]=8'h00; mem['h4CD6]=8'h00; mem['h4CD7]=8'h00;
    mem['h4CD8]=8'h00; mem['h4CD9]=8'h00; mem['h4CDA]=8'h00; mem['h4CDB]=8'h00;
    mem['h4CDC]=8'h00; mem['h4CDD]=8'h00; mem['h4CDE]=8'h00; mem['h4CDF]=8'h00;
    mem['h4CE0]=8'h00; mem['h4CE1]=8'h00; mem['h4CE2]=8'h00; mem['h4CE3]=8'h00;
    mem['h4CE4]=8'h00; mem['h4CE5]=8'h00; mem['h4CE6]=8'h00; mem['h4CE7]=8'h00;
    mem['h4CE8]=8'h00; mem['h4CE9]=8'h00; mem['h4CEA]=8'h00; mem['h4CEB]=8'h00;
    mem['h4CEC]=8'h00; mem['h4CED]=8'h00; mem['h4CEE]=8'h00; mem['h4CEF]=8'h00;
    mem['h4CF0]=8'h00; mem['h4CF1]=8'h00; mem['h4CF2]=8'h00; mem['h4CF3]=8'h00;
    mem['h4CF4]=8'h00; mem['h4CF5]=8'h00; mem['h4CF6]=8'h00; mem['h4CF7]=8'h00;
    mem['h4CF8]=8'h00; mem['h4CF9]=8'h00; mem['h4CFA]=8'h00; mem['h4CFB]=8'h00;
    mem['h4CFC]=8'h00; mem['h4CFD]=8'h00; mem['h4CFE]=8'h00; mem['h4CFF]=8'h00;
    mem['h4D00]=8'h00; mem['h4D01]=8'h00; mem['h4D02]=8'h00; mem['h4D03]=8'h00;
    mem['h4D04]=8'h00; mem['h4D05]=8'h00; mem['h4D06]=8'h00; mem['h4D07]=8'h00;
    mem['h4D08]=8'h00; mem['h4D09]=8'h00; mem['h4D0A]=8'h00; mem['h4D0B]=8'h00;
    mem['h4D0C]=8'h00; mem['h4D0D]=8'h00; mem['h4D0E]=8'h00; mem['h4D0F]=8'h00;
    mem['h4D10]=8'h00; mem['h4D11]=8'h00; mem['h4D12]=8'h00; mem['h4D13]=8'h00;
    mem['h4D14]=8'h00; mem['h4D15]=8'h00; mem['h4D16]=8'h00; mem['h4D17]=8'h00;
    mem['h4D18]=8'h00; mem['h4D19]=8'h00; mem['h4D1A]=8'h00; mem['h4D1B]=8'h00;
    mem['h4D1C]=8'h00; mem['h4D1D]=8'h00; mem['h4D1E]=8'h00; mem['h4D1F]=8'h00;
    mem['h4D20]=8'h00; mem['h4D21]=8'h00; mem['h4D22]=8'h00; mem['h4D23]=8'h00;
    mem['h4D24]=8'h00; mem['h4D25]=8'h00; mem['h4D26]=8'h00; mem['h4D27]=8'h00;
    mem['h4D28]=8'h00; mem['h4D29]=8'h00; mem['h4D2A]=8'h00; mem['h4D2B]=8'h00;
    mem['h4D2C]=8'h00; mem['h4D2D]=8'h00; mem['h4D2E]=8'h00; mem['h4D2F]=8'h00;
    mem['h4D30]=8'h00; mem['h4D31]=8'h00; mem['h4D32]=8'h00; mem['h4D33]=8'h00;
    mem['h4D34]=8'h00; mem['h4D35]=8'h00; mem['h4D36]=8'h00; mem['h4D37]=8'h00;
    mem['h4D38]=8'h00; mem['h4D39]=8'h00; mem['h4D3A]=8'h00; mem['h4D3B]=8'h00;
    mem['h4D3C]=8'h00; mem['h4D3D]=8'h00; mem['h4D3E]=8'h00; mem['h4D3F]=8'h00;
    mem['h4D40]=8'h00; mem['h4D41]=8'h00; mem['h4D42]=8'h00; mem['h4D43]=8'h00;
    mem['h4D44]=8'h00; mem['h4D45]=8'h00; mem['h4D46]=8'h00; mem['h4D47]=8'h00;
    mem['h4D48]=8'h00; mem['h4D49]=8'h00; mem['h4D4A]=8'h00; mem['h4D4B]=8'h00;
    mem['h4D4C]=8'h00; mem['h4D4D]=8'h00; mem['h4D4E]=8'h00; mem['h4D4F]=8'h00;
    mem['h4D50]=8'h00; mem['h4D51]=8'h00; mem['h4D52]=8'h00; mem['h4D53]=8'h00;
    mem['h4D54]=8'h00; mem['h4D55]=8'h00; mem['h4D56]=8'h00; mem['h4D57]=8'h00;
    mem['h4D58]=8'h00; mem['h4D59]=8'h00; mem['h4D5A]=8'h00; mem['h4D5B]=8'h00;
    mem['h4D5C]=8'h00; mem['h4D5D]=8'h00; mem['h4D5E]=8'h00; mem['h4D5F]=8'h00;
    mem['h4D60]=8'h00; mem['h4D61]=8'h00; mem['h4D62]=8'h00; mem['h4D63]=8'h00;
    mem['h4D64]=8'h00; mem['h4D65]=8'h00; mem['h4D66]=8'h00; mem['h4D67]=8'h00;
    mem['h4D68]=8'h00; mem['h4D69]=8'h00; mem['h4D6A]=8'h00; mem['h4D6B]=8'h00;
    mem['h4D6C]=8'h00; mem['h4D6D]=8'h00; mem['h4D6E]=8'h00; mem['h4D6F]=8'h00;
    mem['h4D70]=8'h00; mem['h4D71]=8'h00; mem['h4D72]=8'h00; mem['h4D73]=8'h00;
    mem['h4D74]=8'h00; mem['h4D75]=8'h00; mem['h4D76]=8'h00; mem['h4D77]=8'h00;
    mem['h4D78]=8'h00; mem['h4D79]=8'h00; mem['h4D7A]=8'h00; mem['h4D7B]=8'h00;
    mem['h4D7C]=8'h00; mem['h4D7D]=8'h00; mem['h4D7E]=8'h00; mem['h4D7F]=8'h00;
    mem['h4D80]=8'h00; mem['h4D81]=8'h00; mem['h4D82]=8'h00; mem['h4D83]=8'h00;
    mem['h4D84]=8'h00; mem['h4D85]=8'h00; mem['h4D86]=8'h00; mem['h4D87]=8'h00;
    mem['h4D88]=8'h00; mem['h4D89]=8'h00; mem['h4D8A]=8'h00; mem['h4D8B]=8'h00;
    mem['h4D8C]=8'h00; mem['h4D8D]=8'h00; mem['h4D8E]=8'h00; mem['h4D8F]=8'h00;
    mem['h4D90]=8'h00; mem['h4D91]=8'h00; mem['h4D92]=8'h00; mem['h4D93]=8'h00;
    mem['h4D94]=8'h00; mem['h4D95]=8'h00; mem['h4D96]=8'h00; mem['h4D97]=8'h00;
    mem['h4D98]=8'h00; mem['h4D99]=8'h00; mem['h4D9A]=8'h00; mem['h4D9B]=8'h00;
    mem['h4D9C]=8'h00; mem['h4D9D]=8'h00; mem['h4D9E]=8'h00; mem['h4D9F]=8'h00;
    mem['h4DA0]=8'h00; mem['h4DA1]=8'h00; mem['h4DA2]=8'h00; mem['h4DA3]=8'h00;
    mem['h4DA4]=8'h00; mem['h4DA5]=8'h00; mem['h4DA6]=8'h00; mem['h4DA7]=8'h00;
    mem['h4DA8]=8'h00; mem['h4DA9]=8'h00; mem['h4DAA]=8'h00; mem['h4DAB]=8'h00;
    mem['h4DAC]=8'h00; mem['h4DAD]=8'h00; mem['h4DAE]=8'h00; mem['h4DAF]=8'h00;
    mem['h4DB0]=8'h00; mem['h4DB1]=8'h00; mem['h4DB2]=8'h00; mem['h4DB3]=8'h00;
    mem['h4DB4]=8'h00; mem['h4DB5]=8'h00; mem['h4DB6]=8'h00; mem['h4DB7]=8'h00;
    mem['h4DB8]=8'h00; mem['h4DB9]=8'h00; mem['h4DBA]=8'h00; mem['h4DBB]=8'h00;
    mem['h4DBC]=8'h00; mem['h4DBD]=8'h00; mem['h4DBE]=8'h00; mem['h4DBF]=8'h00;
    mem['h4DC0]=8'h00; mem['h4DC1]=8'h00; mem['h4DC2]=8'h00; mem['h4DC3]=8'h00;
    mem['h4DC4]=8'h00; mem['h4DC5]=8'h00; mem['h4DC6]=8'h00; mem['h4DC7]=8'h00;
    mem['h4DC8]=8'h00; mem['h4DC9]=8'h00; mem['h4DCA]=8'h00; mem['h4DCB]=8'h00;
    mem['h4DCC]=8'h00; mem['h4DCD]=8'h00; mem['h4DCE]=8'h00; mem['h4DCF]=8'h00;
    mem['h4DD0]=8'h00; mem['h4DD1]=8'h00; mem['h4DD2]=8'h00; mem['h4DD3]=8'h00;
    mem['h4DD4]=8'h00; mem['h4DD5]=8'h00; mem['h4DD6]=8'h00; mem['h4DD7]=8'h00;
    mem['h4DD8]=8'h00; mem['h4DD9]=8'h00; mem['h4DDA]=8'h00; mem['h4DDB]=8'h00;
    mem['h4DDC]=8'h00; mem['h4DDD]=8'h00; mem['h4DDE]=8'h00; mem['h4DDF]=8'h00;
    mem['h4DE0]=8'h00; mem['h4DE1]=8'h00; mem['h4DE2]=8'h00; mem['h4DE3]=8'h00;
    mem['h4DE4]=8'h00; mem['h4DE5]=8'h00; mem['h4DE6]=8'h00; mem['h4DE7]=8'h00;
    mem['h4DE8]=8'h00; mem['h4DE9]=8'h00; mem['h4DEA]=8'h00; mem['h4DEB]=8'h00;
    mem['h4DEC]=8'h00; mem['h4DED]=8'h00; mem['h4DEE]=8'h00; mem['h4DEF]=8'h00;
    mem['h4DF0]=8'h00; mem['h4DF1]=8'h00; mem['h4DF2]=8'h00; mem['h4DF3]=8'h00;
    mem['h4DF4]=8'h00; mem['h4DF5]=8'h00; mem['h4DF6]=8'h00; mem['h4DF7]=8'h00;
    mem['h4DF8]=8'h00; mem['h4DF9]=8'h00; mem['h4DFA]=8'h00; mem['h4DFB]=8'h00;
    mem['h4DFC]=8'h00; mem['h4DFD]=8'h00; mem['h4DFE]=8'h00; mem['h4DFF]=8'h00;
    mem['h4E00]=8'h00; mem['h4E01]=8'h00; mem['h4E02]=8'h00; mem['h4E03]=8'h00;
    mem['h4E04]=8'h00; mem['h4E05]=8'h00; mem['h4E06]=8'h00; mem['h4E07]=8'h00;
    mem['h4E08]=8'h00; mem['h4E09]=8'h00; mem['h4E0A]=8'h00; mem['h4E0B]=8'h00;
    mem['h4E0C]=8'h00; mem['h4E0D]=8'h00; mem['h4E0E]=8'h00; mem['h4E0F]=8'h00;
    mem['h4E10]=8'h00; mem['h4E11]=8'h00; mem['h4E12]=8'h00; mem['h4E13]=8'h00;
    mem['h4E14]=8'h00; mem['h4E15]=8'h00; mem['h4E16]=8'h00; mem['h4E17]=8'h00;
    mem['h4E18]=8'h00; mem['h4E19]=8'h00; mem['h4E1A]=8'h00; mem['h4E1B]=8'h00;
    mem['h4E1C]=8'h00; mem['h4E1D]=8'h00; mem['h4E1E]=8'h00; mem['h4E1F]=8'h00;
    mem['h4E20]=8'h00; mem['h4E21]=8'h00; mem['h4E22]=8'h00; mem['h4E23]=8'h00;
    mem['h4E24]=8'h00; mem['h4E25]=8'h00; mem['h4E26]=8'h00; mem['h4E27]=8'h00;
    mem['h4E28]=8'h00; mem['h4E29]=8'h00; mem['h4E2A]=8'h00; mem['h4E2B]=8'h00;
    mem['h4E2C]=8'h00; mem['h4E2D]=8'h00; mem['h4E2E]=8'h00; mem['h4E2F]=8'h00;
    mem['h4E30]=8'h00; mem['h4E31]=8'h00; mem['h4E32]=8'h00; mem['h4E33]=8'h00;
    mem['h4E34]=8'h00; mem['h4E35]=8'h00; mem['h4E36]=8'h00; mem['h4E37]=8'h00;
    mem['h4E38]=8'h00; mem['h4E39]=8'h00; mem['h4E3A]=8'h00; mem['h4E3B]=8'h00;
    mem['h4E3C]=8'h00; mem['h4E3D]=8'h00; mem['h4E3E]=8'h00; mem['h4E3F]=8'h00;
    mem['h4E40]=8'h00; mem['h4E41]=8'h00; mem['h4E42]=8'h00; mem['h4E43]=8'h00;
    mem['h4E44]=8'h00; mem['h4E45]=8'h00; mem['h4E46]=8'h00; mem['h4E47]=8'h00;
    mem['h4E48]=8'h00; mem['h4E49]=8'h00; mem['h4E4A]=8'h00; mem['h4E4B]=8'h00;
    mem['h4E4C]=8'h00; mem['h4E4D]=8'h00; mem['h4E4E]=8'h00; mem['h4E4F]=8'h00;
    mem['h4E50]=8'h00; mem['h4E51]=8'h00; mem['h4E52]=8'h00; mem['h4E53]=8'h00;
    mem['h4E54]=8'h00; mem['h4E55]=8'h00; mem['h4E56]=8'h00; mem['h4E57]=8'h00;
    mem['h4E58]=8'h00; mem['h4E59]=8'h00; mem['h4E5A]=8'h00; mem['h4E5B]=8'h00;
    mem['h4E5C]=8'h00; mem['h4E5D]=8'h00; mem['h4E5E]=8'h00; mem['h4E5F]=8'h00;
    mem['h4E60]=8'h00; mem['h4E61]=8'h00; mem['h4E62]=8'h00; mem['h4E63]=8'h00;
    mem['h4E64]=8'h00; mem['h4E65]=8'h00; mem['h4E66]=8'h00; mem['h4E67]=8'h00;
    mem['h4E68]=8'h00; mem['h4E69]=8'h00; mem['h4E6A]=8'h00; mem['h4E6B]=8'h00;
    mem['h4E6C]=8'h00; mem['h4E6D]=8'h00; mem['h4E6E]=8'h00; mem['h4E6F]=8'h00;
    mem['h4E70]=8'h00; mem['h4E71]=8'h00; mem['h4E72]=8'h00; mem['h4E73]=8'h00;
    mem['h4E74]=8'h00; mem['h4E75]=8'h00; mem['h4E76]=8'h00; mem['h4E77]=8'h00;
    mem['h4E78]=8'h00; mem['h4E79]=8'h00; mem['h4E7A]=8'h00; mem['h4E7B]=8'h00;
    mem['h4E7C]=8'h00; mem['h4E7D]=8'h00; mem['h4E7E]=8'h00; mem['h4E7F]=8'h00;
    mem['h4E80]=8'h00; mem['h4E81]=8'h00; mem['h4E82]=8'h00; mem['h4E83]=8'h00;
    mem['h4E84]=8'h00; mem['h4E85]=8'h00; mem['h4E86]=8'h00; mem['h4E87]=8'h00;
    mem['h4E88]=8'h00; mem['h4E89]=8'h00; mem['h4E8A]=8'h00; mem['h4E8B]=8'h00;
    mem['h4E8C]=8'h00; mem['h4E8D]=8'h00; mem['h4E8E]=8'h00; mem['h4E8F]=8'h00;
    mem['h4E90]=8'h00; mem['h4E91]=8'h00; mem['h4E92]=8'h00; mem['h4E93]=8'h00;
    mem['h4E94]=8'h00; mem['h4E95]=8'h00; mem['h4E96]=8'h00; mem['h4E97]=8'h00;
    mem['h4E98]=8'h00; mem['h4E99]=8'h00; mem['h4E9A]=8'h00; mem['h4E9B]=8'h00;
    mem['h4E9C]=8'h00; mem['h4E9D]=8'h00; mem['h4E9E]=8'h00; mem['h4E9F]=8'h00;
    mem['h4EA0]=8'h00; mem['h4EA1]=8'h00; mem['h4EA2]=8'h00; mem['h4EA3]=8'h00;
    mem['h4EA4]=8'h00; mem['h4EA5]=8'h00; mem['h4EA6]=8'h00; mem['h4EA7]=8'h00;
    mem['h4EA8]=8'h00; mem['h4EA9]=8'h00; mem['h4EAA]=8'h00; mem['h4EAB]=8'h00;
    mem['h4EAC]=8'h00; mem['h4EAD]=8'h00; mem['h4EAE]=8'h00; mem['h4EAF]=8'h00;
    mem['h4EB0]=8'h00; mem['h4EB1]=8'h00; mem['h4EB2]=8'h00; mem['h4EB3]=8'h00;
    mem['h4EB4]=8'h00; mem['h4EB5]=8'h00; mem['h4EB6]=8'h00; mem['h4EB7]=8'h00;
    mem['h4EB8]=8'h00; mem['h4EB9]=8'h00; mem['h4EBA]=8'h00; mem['h4EBB]=8'h00;
    mem['h4EBC]=8'h00; mem['h4EBD]=8'h00; mem['h4EBE]=8'h00; mem['h4EBF]=8'h00;
    mem['h4EC0]=8'h00; mem['h4EC1]=8'h00; mem['h4EC2]=8'h00; mem['h4EC3]=8'h00;
    mem['h4EC4]=8'h00; mem['h4EC5]=8'h00; mem['h4EC6]=8'h00; mem['h4EC7]=8'h00;
    mem['h4EC8]=8'h00; mem['h4EC9]=8'h00; mem['h4ECA]=8'h00; mem['h4ECB]=8'h00;
    mem['h4ECC]=8'h00; mem['h4ECD]=8'h00; mem['h4ECE]=8'h00; mem['h4ECF]=8'h00;
    mem['h4ED0]=8'h00; mem['h4ED1]=8'h00; mem['h4ED2]=8'h00; mem['h4ED3]=8'h00;
    mem['h4ED4]=8'h00; mem['h4ED5]=8'h00; mem['h4ED6]=8'h00; mem['h4ED7]=8'h00;
    mem['h4ED8]=8'h00; mem['h4ED9]=8'h00; mem['h4EDA]=8'h00; mem['h4EDB]=8'h00;
    mem['h4EDC]=8'h00; mem['h4EDD]=8'h00; mem['h4EDE]=8'h00; mem['h4EDF]=8'h00;
    mem['h4EE0]=8'h00; mem['h4EE1]=8'h00; mem['h4EE2]=8'h00; mem['h4EE3]=8'h00;
    mem['h4EE4]=8'h00; mem['h4EE5]=8'h00; mem['h4EE6]=8'h00; mem['h4EE7]=8'h00;
    mem['h4EE8]=8'h00; mem['h4EE9]=8'h00; mem['h4EEA]=8'h00; mem['h4EEB]=8'h00;
    mem['h4EEC]=8'h00; mem['h4EED]=8'h00; mem['h4EEE]=8'h00; mem['h4EEF]=8'h00;
    mem['h4EF0]=8'h00; mem['h4EF1]=8'h00; mem['h4EF2]=8'h00; mem['h4EF3]=8'h00;
    mem['h4EF4]=8'h00; mem['h4EF5]=8'h00; mem['h4EF6]=8'h00; mem['h4EF7]=8'h00;
    mem['h4EF8]=8'h00; mem['h4EF9]=8'h00; mem['h4EFA]=8'h00; mem['h4EFB]=8'h00;
    mem['h4EFC]=8'h00; mem['h4EFD]=8'h00; mem['h4EFE]=8'h00; mem['h4EFF]=8'h00;
    mem['h4F00]=8'h00; mem['h4F01]=8'h00; mem['h4F02]=8'h00; mem['h4F03]=8'h00;
    mem['h4F04]=8'h00; mem['h4F05]=8'h00; mem['h4F06]=8'h00; mem['h4F07]=8'h00;
    mem['h4F08]=8'h00; mem['h4F09]=8'h00; mem['h4F0A]=8'h00; mem['h4F0B]=8'h00;
    mem['h4F0C]=8'h00; mem['h4F0D]=8'h00; mem['h4F0E]=8'h00; mem['h4F0F]=8'h00;
    mem['h4F10]=8'h00; mem['h4F11]=8'h00; mem['h4F12]=8'h00; mem['h4F13]=8'h00;
    mem['h4F14]=8'h00; mem['h4F15]=8'h00; mem['h4F16]=8'h00; mem['h4F17]=8'h00;
    mem['h4F18]=8'h00; mem['h4F19]=8'h00; mem['h4F1A]=8'h00; mem['h4F1B]=8'h00;
    mem['h4F1C]=8'h00; mem['h4F1D]=8'h00; mem['h4F1E]=8'h00; mem['h4F1F]=8'h00;
    mem['h4F20]=8'h00; mem['h4F21]=8'h00; mem['h4F22]=8'h00; mem['h4F23]=8'h00;
    mem['h4F24]=8'h00; mem['h4F25]=8'h00; mem['h4F26]=8'h00; mem['h4F27]=8'h00;
    mem['h4F28]=8'h00; mem['h4F29]=8'h00; mem['h4F2A]=8'h00; mem['h4F2B]=8'h00;
    mem['h4F2C]=8'h00; mem['h4F2D]=8'h00; mem['h4F2E]=8'h00; mem['h4F2F]=8'h00;
    mem['h4F30]=8'h00; mem['h4F31]=8'h00; mem['h4F32]=8'h00; mem['h4F33]=8'h00;
    mem['h4F34]=8'h00; mem['h4F35]=8'h00; mem['h4F36]=8'h00; mem['h4F37]=8'h00;
    mem['h4F38]=8'h00; mem['h4F39]=8'h00; mem['h4F3A]=8'h00; mem['h4F3B]=8'h00;
    mem['h4F3C]=8'h00; mem['h4F3D]=8'h00; mem['h4F3E]=8'h00; mem['h4F3F]=8'h00;
    mem['h4F40]=8'h00; mem['h4F41]=8'h00; mem['h4F42]=8'h00; mem['h4F43]=8'h00;
    mem['h4F44]=8'h00; mem['h4F45]=8'h00; mem['h4F46]=8'h00; mem['h4F47]=8'h00;
    mem['h4F48]=8'h00; mem['h4F49]=8'h00; mem['h4F4A]=8'h00; mem['h4F4B]=8'h00;
    mem['h4F4C]=8'h00; mem['h4F4D]=8'h00; mem['h4F4E]=8'h00; mem['h4F4F]=8'h00;
    mem['h4F50]=8'h00; mem['h4F51]=8'h00; mem['h4F52]=8'h00; mem['h4F53]=8'h00;
    mem['h4F54]=8'h00; mem['h4F55]=8'h00; mem['h4F56]=8'h00; mem['h4F57]=8'h00;
    mem['h4F58]=8'h00; mem['h4F59]=8'h00; mem['h4F5A]=8'h00; mem['h4F5B]=8'h00;
    mem['h4F5C]=8'h00; mem['h4F5D]=8'h00; mem['h4F5E]=8'h00; mem['h4F5F]=8'h00;
    mem['h4F60]=8'h00; mem['h4F61]=8'h00; mem['h4F62]=8'h00; mem['h4F63]=8'h00;
    mem['h4F64]=8'h00; mem['h4F65]=8'h00; mem['h4F66]=8'h00; mem['h4F67]=8'h00;
    mem['h4F68]=8'h00; mem['h4F69]=8'h00; mem['h4F6A]=8'h00; mem['h4F6B]=8'h00;
    mem['h4F6C]=8'h00; mem['h4F6D]=8'h00; mem['h4F6E]=8'h00; mem['h4F6F]=8'h00;
    mem['h4F70]=8'h00; mem['h4F71]=8'h00; mem['h4F72]=8'h00; mem['h4F73]=8'h00;
    mem['h4F74]=8'h00; mem['h4F75]=8'h00; mem['h4F76]=8'h00; mem['h4F77]=8'h00;
    mem['h4F78]=8'h00; mem['h4F79]=8'h00; mem['h4F7A]=8'h00; mem['h4F7B]=8'h00;
    mem['h4F7C]=8'h00; mem['h4F7D]=8'h00; mem['h4F7E]=8'h00; mem['h4F7F]=8'h00;
    mem['h4F80]=8'h00; mem['h4F81]=8'h00; mem['h4F82]=8'h00; mem['h4F83]=8'h00;
    mem['h4F84]=8'h00; mem['h4F85]=8'h00; mem['h4F86]=8'h00; mem['h4F87]=8'h00;
    mem['h4F88]=8'h00; mem['h4F89]=8'h00; mem['h4F8A]=8'h00; mem['h4F8B]=8'h00;
    mem['h4F8C]=8'h00; mem['h4F8D]=8'h00; mem['h4F8E]=8'h00; mem['h4F8F]=8'h00;
    mem['h4F90]=8'h00; mem['h4F91]=8'h00; mem['h4F92]=8'h00; mem['h4F93]=8'h00;
    mem['h4F94]=8'h00; mem['h4F95]=8'h00; mem['h4F96]=8'h00; mem['h4F97]=8'h00;
    mem['h4F98]=8'h00; mem['h4F99]=8'h00; mem['h4F9A]=8'h00; mem['h4F9B]=8'h00;
    mem['h4F9C]=8'h00; mem['h4F9D]=8'h00; mem['h4F9E]=8'h00; mem['h4F9F]=8'h00;
    mem['h4FA0]=8'h00; mem['h4FA1]=8'h00; mem['h4FA2]=8'h00; mem['h4FA3]=8'h00;
    mem['h4FA4]=8'h00; mem['h4FA5]=8'h00; mem['h4FA6]=8'h00; mem['h4FA7]=8'h00;
    mem['h4FA8]=8'h00; mem['h4FA9]=8'h00; mem['h4FAA]=8'h00; mem['h4FAB]=8'h00;
    mem['h4FAC]=8'h00; mem['h4FAD]=8'h00; mem['h4FAE]=8'h00; mem['h4FAF]=8'h00;
    mem['h4FB0]=8'h00; mem['h4FB1]=8'h00; mem['h4FB2]=8'h00; mem['h4FB3]=8'h00;
    mem['h4FB4]=8'h00; mem['h4FB5]=8'h00; mem['h4FB6]=8'h00; mem['h4FB7]=8'h00;
    mem['h4FB8]=8'h00; mem['h4FB9]=8'h00; mem['h4FBA]=8'h00; mem['h4FBB]=8'h00;
    mem['h4FBC]=8'h00; mem['h4FBD]=8'h00; mem['h4FBE]=8'h00; mem['h4FBF]=8'h00;
    mem['h4FC0]=8'h00; mem['h4FC1]=8'h00; mem['h4FC2]=8'h00; mem['h4FC3]=8'h00;
    mem['h4FC4]=8'h00; mem['h4FC5]=8'h00; mem['h4FC6]=8'h00; mem['h4FC7]=8'h00;
    mem['h4FC8]=8'h00; mem['h4FC9]=8'h00; mem['h4FCA]=8'h00; mem['h4FCB]=8'h00;
    mem['h4FCC]=8'h00; mem['h4FCD]=8'h00; mem['h4FCE]=8'h00; mem['h4FCF]=8'h00;
    mem['h4FD0]=8'h00; mem['h4FD1]=8'h00; mem['h4FD2]=8'h00; mem['h4FD3]=8'h00;
    mem['h4FD4]=8'h00; mem['h4FD5]=8'h00; mem['h4FD6]=8'h00; mem['h4FD7]=8'h00;
    mem['h4FD8]=8'h00; mem['h4FD9]=8'h00; mem['h4FDA]=8'h00; mem['h4FDB]=8'h00;
    mem['h4FDC]=8'h00; mem['h4FDD]=8'h00; mem['h4FDE]=8'h00; mem['h4FDF]=8'h00;
    mem['h4FE0]=8'h00; mem['h4FE1]=8'h00; mem['h4FE2]=8'h00; mem['h4FE3]=8'h00;
    mem['h4FE4]=8'h00; mem['h4FE5]=8'h00; mem['h4FE6]=8'h00; mem['h4FE7]=8'h00;
    mem['h4FE8]=8'h00; mem['h4FE9]=8'h00; mem['h4FEA]=8'h00; mem['h4FEB]=8'h00;
    mem['h4FEC]=8'h00; mem['h4FED]=8'h00; mem['h4FEE]=8'h00; mem['h4FEF]=8'h00;
    mem['h4FF0]=8'h00; mem['h4FF1]=8'h00; mem['h4FF2]=8'h00; mem['h4FF3]=8'h00;
    mem['h4FF4]=8'h00; mem['h4FF5]=8'h00; mem['h4FF6]=8'h00; mem['h4FF7]=8'h00;
    mem['h4FF8]=8'h00; mem['h4FF9]=8'h00; mem['h4FFA]=8'h00; mem['h4FFB]=8'h00;
    mem['h4FFC]=8'h00; mem['h4FFD]=8'h00; mem['h4FFE]=8'h00; mem['h4FFF]=8'h00;
    mem['h5000]=8'h00; mem['h5001]=8'h00; mem['h5002]=8'h00; mem['h5003]=8'h00;
    mem['h5004]=8'h00; mem['h5005]=8'h00; mem['h5006]=8'h00; mem['h5007]=8'h00;
    mem['h5008]=8'h00; mem['h5009]=8'h00; mem['h500A]=8'h00; mem['h500B]=8'h00;
    mem['h500C]=8'h00; mem['h500D]=8'h00; mem['h500E]=8'h00; mem['h500F]=8'h00;
    mem['h5010]=8'h00; mem['h5011]=8'h00; mem['h5012]=8'h00; mem['h5013]=8'h00;
    mem['h5014]=8'h00; mem['h5015]=8'h00; mem['h5016]=8'h00; mem['h5017]=8'h00;
    mem['h5018]=8'h00; mem['h5019]=8'h00; mem['h501A]=8'h00; mem['h501B]=8'h00;
    mem['h501C]=8'h00; mem['h501D]=8'h00; mem['h501E]=8'h00; mem['h501F]=8'h00;
    mem['h5020]=8'h00; mem['h5021]=8'h00; mem['h5022]=8'h00; mem['h5023]=8'h00;
    mem['h5024]=8'h00; mem['h5025]=8'h00; mem['h5026]=8'h00; mem['h5027]=8'h00;
    mem['h5028]=8'h00; mem['h5029]=8'h00; mem['h502A]=8'h00; mem['h502B]=8'h00;
    mem['h502C]=8'h00; mem['h502D]=8'h00; mem['h502E]=8'h00; mem['h502F]=8'h00;
    mem['h5030]=8'h00; mem['h5031]=8'h00; mem['h5032]=8'h00; mem['h5033]=8'h00;
    mem['h5034]=8'h00; mem['h5035]=8'h00; mem['h5036]=8'h00; mem['h5037]=8'h00;
    mem['h5038]=8'h00; mem['h5039]=8'h00; mem['h503A]=8'h00; mem['h503B]=8'h00;
    mem['h503C]=8'h00; mem['h503D]=8'h00; mem['h503E]=8'h00; mem['h503F]=8'h00;
    mem['h5040]=8'h00; mem['h5041]=8'h00; mem['h5042]=8'h00; mem['h5043]=8'h00;
    mem['h5044]=8'h00; mem['h5045]=8'h00; mem['h5046]=8'h00; mem['h5047]=8'h00;
    mem['h5048]=8'h00; mem['h5049]=8'h00; mem['h504A]=8'h00; mem['h504B]=8'h00;
    mem['h504C]=8'h00; mem['h504D]=8'h00; mem['h504E]=8'h00; mem['h504F]=8'h00;
    mem['h5050]=8'h00; mem['h5051]=8'h00; mem['h5052]=8'h00; mem['h5053]=8'h00;
    mem['h5054]=8'h00; mem['h5055]=8'h00; mem['h5056]=8'h00; mem['h5057]=8'h00;
    mem['h5058]=8'h00; mem['h5059]=8'h00; mem['h505A]=8'h00; mem['h505B]=8'h00;
    mem['h505C]=8'h00; mem['h505D]=8'h00; mem['h505E]=8'h00; mem['h505F]=8'h00;
    mem['h5060]=8'h00; mem['h5061]=8'h00; mem['h5062]=8'h00; mem['h5063]=8'h00;
    mem['h5064]=8'h00; mem['h5065]=8'h00; mem['h5066]=8'h00; mem['h5067]=8'h00;
    mem['h5068]=8'h00; mem['h5069]=8'h00; mem['h506A]=8'h00; mem['h506B]=8'h00;
    mem['h506C]=8'h00; mem['h506D]=8'h00; mem['h506E]=8'h00; mem['h506F]=8'h00;
    mem['h5070]=8'h00; mem['h5071]=8'h00; mem['h5072]=8'h00; mem['h5073]=8'h00;
    mem['h5074]=8'h00; mem['h5075]=8'h00; mem['h5076]=8'h00; mem['h5077]=8'h00;
    mem['h5078]=8'h00; mem['h5079]=8'h00; mem['h507A]=8'h00; mem['h507B]=8'h00;
    mem['h507C]=8'h00; mem['h507D]=8'h00; mem['h507E]=8'h00; mem['h507F]=8'h00;
    mem['h5080]=8'h00; mem['h5081]=8'h00; mem['h5082]=8'h00; mem['h5083]=8'h00;
    mem['h5084]=8'h00; mem['h5085]=8'h00; mem['h5086]=8'h00; mem['h5087]=8'h00;
    mem['h5088]=8'h00; mem['h5089]=8'h00; mem['h508A]=8'h00; mem['h508B]=8'h00;
    mem['h508C]=8'h00; mem['h508D]=8'h00; mem['h508E]=8'h00; mem['h508F]=8'h00;
    mem['h5090]=8'h00; mem['h5091]=8'h00; mem['h5092]=8'h00; mem['h5093]=8'h00;
    mem['h5094]=8'h00; mem['h5095]=8'h00; mem['h5096]=8'h00; mem['h5097]=8'h00;
    mem['h5098]=8'h00; mem['h5099]=8'h00; mem['h509A]=8'h00; mem['h509B]=8'h00;
    mem['h509C]=8'h00; mem['h509D]=8'h00; mem['h509E]=8'h00; mem['h509F]=8'h00;
    mem['h50A0]=8'h00; mem['h50A1]=8'h00; mem['h50A2]=8'h00; mem['h50A3]=8'h00;
    mem['h50A4]=8'h00; mem['h50A5]=8'h00; mem['h50A6]=8'h00; mem['h50A7]=8'h00;
    mem['h50A8]=8'h00; mem['h50A9]=8'h00; mem['h50AA]=8'h00; mem['h50AB]=8'h00;
    mem['h50AC]=8'h00; mem['h50AD]=8'h00; mem['h50AE]=8'h00; mem['h50AF]=8'h00;
    mem['h50B0]=8'h00; mem['h50B1]=8'h00; mem['h50B2]=8'h00; mem['h50B3]=8'h00;
    mem['h50B4]=8'h00; mem['h50B5]=8'h00; mem['h50B6]=8'h00; mem['h50B7]=8'h00;
    mem['h50B8]=8'h00; mem['h50B9]=8'h00; mem['h50BA]=8'h00; mem['h50BB]=8'h00;
    mem['h50BC]=8'h00; mem['h50BD]=8'h00; mem['h50BE]=8'h00; mem['h50BF]=8'h00;
    mem['h50C0]=8'h00; mem['h50C1]=8'h00; mem['h50C2]=8'h00; mem['h50C3]=8'h00;
    mem['h50C4]=8'h00; mem['h50C5]=8'h00; mem['h50C6]=8'h00; mem['h50C7]=8'h00;
    mem['h50C8]=8'h00; mem['h50C9]=8'h00; mem['h50CA]=8'h00; mem['h50CB]=8'h00;
    mem['h50CC]=8'h00; mem['h50CD]=8'h00; mem['h50CE]=8'h00; mem['h50CF]=8'h00;
    mem['h50D0]=8'h00; mem['h50D1]=8'h00; mem['h50D2]=8'h00; mem['h50D3]=8'h00;
    mem['h50D4]=8'h00; mem['h50D5]=8'h00; mem['h50D6]=8'h00; mem['h50D7]=8'h00;
    mem['h50D8]=8'h00; mem['h50D9]=8'h00; mem['h50DA]=8'h00; mem['h50DB]=8'h00;
    mem['h50DC]=8'h00; mem['h50DD]=8'h00; mem['h50DE]=8'h00; mem['h50DF]=8'h00;
    mem['h50E0]=8'h00; mem['h50E1]=8'h00; mem['h50E2]=8'h00; mem['h50E3]=8'h00;
    mem['h50E4]=8'h00; mem['h50E5]=8'h00; mem['h50E6]=8'h00; mem['h50E7]=8'h00;
    mem['h50E8]=8'h00; mem['h50E9]=8'h00; mem['h50EA]=8'h00; mem['h50EB]=8'h00;
    mem['h50EC]=8'h00; mem['h50ED]=8'h00; mem['h50EE]=8'h00; mem['h50EF]=8'h00;
    mem['h50F0]=8'h00; mem['h50F1]=8'h00; mem['h50F2]=8'h00; mem['h50F3]=8'h00;
    mem['h50F4]=8'h00; mem['h50F5]=8'h00; mem['h50F6]=8'h00; mem['h50F7]=8'h00;
    mem['h50F8]=8'h00; mem['h50F9]=8'h00; mem['h50FA]=8'h00; mem['h50FB]=8'h00;
    mem['h50FC]=8'h00; mem['h50FD]=8'h00; mem['h50FE]=8'h00; mem['h50FF]=8'h00;
    mem['h5100]=8'h00; mem['h5101]=8'h00; mem['h5102]=8'h00; mem['h5103]=8'h00;
    mem['h5104]=8'h00; mem['h5105]=8'h00; mem['h5106]=8'h00; mem['h5107]=8'h00;
    mem['h5108]=8'h00; mem['h5109]=8'h00; mem['h510A]=8'h00; mem['h510B]=8'h00;
    mem['h510C]=8'h00; mem['h510D]=8'h00; mem['h510E]=8'h00; mem['h510F]=8'h00;
    mem['h5110]=8'h00; mem['h5111]=8'h00; mem['h5112]=8'h00; mem['h5113]=8'h00;
    mem['h5114]=8'h00; mem['h5115]=8'h00; mem['h5116]=8'h00; mem['h5117]=8'h00;
    mem['h5118]=8'h00; mem['h5119]=8'h00; mem['h511A]=8'h00; mem['h511B]=8'h00;
    mem['h511C]=8'h00; mem['h511D]=8'h00; mem['h511E]=8'h00; mem['h511F]=8'h00;
    mem['h5120]=8'h00; mem['h5121]=8'h00; mem['h5122]=8'h00; mem['h5123]=8'h00;
    mem['h5124]=8'h00; mem['h5125]=8'h00; mem['h5126]=8'h00; mem['h5127]=8'h00;
    mem['h5128]=8'h00; mem['h5129]=8'h00; mem['h512A]=8'h00; mem['h512B]=8'h00;
    mem['h512C]=8'h00; mem['h512D]=8'h00; mem['h512E]=8'h00; mem['h512F]=8'h00;
    mem['h5130]=8'h00; mem['h5131]=8'h00; mem['h5132]=8'h00; mem['h5133]=8'h00;
    mem['h5134]=8'h00; mem['h5135]=8'h00; mem['h5136]=8'h00; mem['h5137]=8'h00;
    mem['h5138]=8'h00; mem['h5139]=8'h00; mem['h513A]=8'h00; mem['h513B]=8'h00;
    mem['h513C]=8'h00; mem['h513D]=8'h00; mem['h513E]=8'h00; mem['h513F]=8'h00;
    mem['h5140]=8'h00; mem['h5141]=8'h00; mem['h5142]=8'h00; mem['h5143]=8'h00;
    mem['h5144]=8'h00; mem['h5145]=8'h00; mem['h5146]=8'h00; mem['h5147]=8'h00;
    mem['h5148]=8'h00; mem['h5149]=8'h00; mem['h514A]=8'h00; mem['h514B]=8'h00;
    mem['h514C]=8'h00; mem['h514D]=8'h00; mem['h514E]=8'h00; mem['h514F]=8'h00;
    mem['h5150]=8'h00; mem['h5151]=8'h00; mem['h5152]=8'h00; mem['h5153]=8'h00;
    mem['h5154]=8'h00; mem['h5155]=8'h00; mem['h5156]=8'h00; mem['h5157]=8'h00;
    mem['h5158]=8'h00; mem['h5159]=8'h00; mem['h515A]=8'h00; mem['h515B]=8'h00;
    mem['h515C]=8'h00; mem['h515D]=8'h00; mem['h515E]=8'h00; mem['h515F]=8'h00;
    mem['h5160]=8'h00; mem['h5161]=8'h00; mem['h5162]=8'h00; mem['h5163]=8'h00;
    mem['h5164]=8'h00; mem['h5165]=8'h00; mem['h5166]=8'h00; mem['h5167]=8'h00;
    mem['h5168]=8'h00; mem['h5169]=8'h00; mem['h516A]=8'h00; mem['h516B]=8'h00;
    mem['h516C]=8'h00; mem['h516D]=8'h00; mem['h516E]=8'h00; mem['h516F]=8'h00;
    mem['h5170]=8'h00; mem['h5171]=8'h00; mem['h5172]=8'h00; mem['h5173]=8'h00;
    mem['h5174]=8'h00; mem['h5175]=8'h00; mem['h5176]=8'h00; mem['h5177]=8'h00;
    mem['h5178]=8'h00; mem['h5179]=8'h00; mem['h517A]=8'h00; mem['h517B]=8'h00;
    mem['h517C]=8'h00; mem['h517D]=8'h00; mem['h517E]=8'h00; mem['h517F]=8'h00;
    mem['h5180]=8'h00; mem['h5181]=8'h00; mem['h5182]=8'h00; mem['h5183]=8'h00;
    mem['h5184]=8'h00; mem['h5185]=8'h00; mem['h5186]=8'h00; mem['h5187]=8'h00;
    mem['h5188]=8'h00; mem['h5189]=8'h00; mem['h518A]=8'h00; mem['h518B]=8'h00;
    mem['h518C]=8'h00; mem['h518D]=8'h00; mem['h518E]=8'h00; mem['h518F]=8'h00;
    mem['h5190]=8'h00; mem['h5191]=8'h00; mem['h5192]=8'h00; mem['h5193]=8'h00;
    mem['h5194]=8'h00; mem['h5195]=8'h00; mem['h5196]=8'h00; mem['h5197]=8'h00;
    mem['h5198]=8'h00; mem['h5199]=8'h00; mem['h519A]=8'h00; mem['h519B]=8'h00;
    mem['h519C]=8'h00; mem['h519D]=8'h00; mem['h519E]=8'h00; mem['h519F]=8'h00;
    mem['h51A0]=8'h00; mem['h51A1]=8'h00; mem['h51A2]=8'h00; mem['h51A3]=8'h00;
    mem['h51A4]=8'h00; mem['h51A5]=8'h00; mem['h51A6]=8'h00; mem['h51A7]=8'h00;
    mem['h51A8]=8'h00; mem['h51A9]=8'h00; mem['h51AA]=8'h00; mem['h51AB]=8'h00;
    mem['h51AC]=8'h00; mem['h51AD]=8'h00; mem['h51AE]=8'h00; mem['h51AF]=8'h00;
    mem['h51B0]=8'h00; mem['h51B1]=8'h00; mem['h51B2]=8'h00; mem['h51B3]=8'h00;
    mem['h51B4]=8'h00; mem['h51B5]=8'h00; mem['h51B6]=8'h00; mem['h51B7]=8'h00;
    mem['h51B8]=8'h00; mem['h51B9]=8'h00; mem['h51BA]=8'h00; mem['h51BB]=8'h00;
    mem['h51BC]=8'h00; mem['h51BD]=8'h00; mem['h51BE]=8'h00; mem['h51BF]=8'h00;
    mem['h51C0]=8'h00; mem['h51C1]=8'h00; mem['h51C2]=8'h00; mem['h51C3]=8'h00;
    mem['h51C4]=8'h00; mem['h51C5]=8'h00; mem['h51C6]=8'h00; mem['h51C7]=8'h00;
    mem['h51C8]=8'h00; mem['h51C9]=8'h00; mem['h51CA]=8'h00; mem['h51CB]=8'h00;
    mem['h51CC]=8'h00; mem['h51CD]=8'h00; mem['h51CE]=8'h00; mem['h51CF]=8'h00;
    mem['h51D0]=8'h00; mem['h51D1]=8'h00; mem['h51D2]=8'h00; mem['h51D3]=8'h00;
    mem['h51D4]=8'h00; mem['h51D5]=8'h00; mem['h51D6]=8'h00; mem['h51D7]=8'h00;
    mem['h51D8]=8'h00; mem['h51D9]=8'h00; mem['h51DA]=8'h00; mem['h51DB]=8'h00;
    mem['h51DC]=8'h00; mem['h51DD]=8'h00; mem['h51DE]=8'h00; mem['h51DF]=8'h00;
    mem['h51E0]=8'h00; mem['h51E1]=8'h00; mem['h51E2]=8'h00; mem['h51E3]=8'h00;
    mem['h51E4]=8'h00; mem['h51E5]=8'h00; mem['h51E6]=8'h00; mem['h51E7]=8'h00;
    mem['h51E8]=8'h00; mem['h51E9]=8'h00; mem['h51EA]=8'h00; mem['h51EB]=8'h00;
    mem['h51EC]=8'h00; mem['h51ED]=8'h00; mem['h51EE]=8'h00; mem['h51EF]=8'h00;
    mem['h51F0]=8'h00; mem['h51F1]=8'h00; mem['h51F2]=8'h00; mem['h51F3]=8'h00;
    mem['h51F4]=8'h00; mem['h51F5]=8'h00; mem['h51F6]=8'h00; mem['h51F7]=8'h00;
    mem['h51F8]=8'h00; mem['h51F9]=8'h00; mem['h51FA]=8'h00; mem['h51FB]=8'h00;
    mem['h51FC]=8'h00; mem['h51FD]=8'h00; mem['h51FE]=8'h00; mem['h51FF]=8'h00;
    mem['h5200]=8'h00; mem['h5201]=8'h00; mem['h5202]=8'h00; mem['h5203]=8'h00;
    mem['h5204]=8'h00; mem['h5205]=8'h00; mem['h5206]=8'h00; mem['h5207]=8'h00;
    mem['h5208]=8'h00; mem['h5209]=8'h00; mem['h520A]=8'h00; mem['h520B]=8'h00;
    mem['h520C]=8'h00; mem['h520D]=8'h00; mem['h520E]=8'h00; mem['h520F]=8'h00;
    mem['h5210]=8'h00; mem['h5211]=8'h00; mem['h5212]=8'h00; mem['h5213]=8'h00;
    mem['h5214]=8'h00; mem['h5215]=8'h00; mem['h5216]=8'h00; mem['h5217]=8'h00;
    mem['h5218]=8'h00; mem['h5219]=8'h00; mem['h521A]=8'h00; mem['h521B]=8'h00;
    mem['h521C]=8'h00; mem['h521D]=8'h00; mem['h521E]=8'h00; mem['h521F]=8'h00;
    mem['h5220]=8'h00; mem['h5221]=8'h00; mem['h5222]=8'h00; mem['h5223]=8'h00;
    mem['h5224]=8'h00; mem['h5225]=8'h00; mem['h5226]=8'h00; mem['h5227]=8'h00;
    mem['h5228]=8'h00; mem['h5229]=8'h00; mem['h522A]=8'h00; mem['h522B]=8'h00;
    mem['h522C]=8'h00; mem['h522D]=8'h00; mem['h522E]=8'h00; mem['h522F]=8'h00;
    mem['h5230]=8'h00; mem['h5231]=8'h00; mem['h5232]=8'h00; mem['h5233]=8'h00;
    mem['h5234]=8'h00; mem['h5235]=8'h00; mem['h5236]=8'h00; mem['h5237]=8'h00;
    mem['h5238]=8'h00; mem['h5239]=8'h00; mem['h523A]=8'h00; mem['h523B]=8'h00;
    mem['h523C]=8'h00; mem['h523D]=8'h00; mem['h523E]=8'h00; mem['h523F]=8'h00;
    mem['h5240]=8'h00; mem['h5241]=8'h00; mem['h5242]=8'h00; mem['h5243]=8'h00;
    mem['h5244]=8'h00; mem['h5245]=8'h00; mem['h5246]=8'h00; mem['h5247]=8'h00;
    mem['h5248]=8'h00; mem['h5249]=8'h00; mem['h524A]=8'h00; mem['h524B]=8'h00;
    mem['h524C]=8'h00; mem['h524D]=8'h00; mem['h524E]=8'h00; mem['h524F]=8'h00;
    mem['h5250]=8'h00; mem['h5251]=8'h00; mem['h5252]=8'h00; mem['h5253]=8'h00;
    mem['h5254]=8'h00; mem['h5255]=8'h00; mem['h5256]=8'h00; mem['h5257]=8'h00;
    mem['h5258]=8'h00; mem['h5259]=8'h00; mem['h525A]=8'h00; mem['h525B]=8'h00;
    mem['h525C]=8'h00; mem['h525D]=8'h00; mem['h525E]=8'h00; mem['h525F]=8'h00;
    mem['h5260]=8'h00; mem['h5261]=8'h00; mem['h5262]=8'h00; mem['h5263]=8'h00;
    mem['h5264]=8'h00; mem['h5265]=8'h00; mem['h5266]=8'h00; mem['h5267]=8'h00;
    mem['h5268]=8'h00; mem['h5269]=8'h00; mem['h526A]=8'h00; mem['h526B]=8'h00;
    mem['h526C]=8'h00; mem['h526D]=8'h00; mem['h526E]=8'h00; mem['h526F]=8'h00;
    mem['h5270]=8'h00; mem['h5271]=8'h00; mem['h5272]=8'h00; mem['h5273]=8'h00;
    mem['h5274]=8'h00; mem['h5275]=8'h00; mem['h5276]=8'h00; mem['h5277]=8'h00;
    mem['h5278]=8'h00; mem['h5279]=8'h00; mem['h527A]=8'h00; mem['h527B]=8'h00;
    mem['h527C]=8'h00; mem['h527D]=8'h00; mem['h527E]=8'h00; mem['h527F]=8'h00;
    mem['h5280]=8'h00; mem['h5281]=8'h00; mem['h5282]=8'h00; mem['h5283]=8'h00;
    mem['h5284]=8'h00; mem['h5285]=8'h00; mem['h5286]=8'h00; mem['h5287]=8'h00;
    mem['h5288]=8'h00; mem['h5289]=8'h00; mem['h528A]=8'h00; mem['h528B]=8'h00;
    mem['h528C]=8'h00; mem['h528D]=8'h00; mem['h528E]=8'h00; mem['h528F]=8'h00;
    mem['h5290]=8'h00; mem['h5291]=8'h00; mem['h5292]=8'h00; mem['h5293]=8'h00;
    mem['h5294]=8'h00; mem['h5295]=8'h00; mem['h5296]=8'h00; mem['h5297]=8'h00;
    mem['h5298]=8'h00; mem['h5299]=8'h00; mem['h529A]=8'h00; mem['h529B]=8'h00;
    mem['h529C]=8'h00; mem['h529D]=8'h00; mem['h529E]=8'h00; mem['h529F]=8'h00;
    mem['h52A0]=8'h00; mem['h52A1]=8'h00; mem['h52A2]=8'h00; mem['h52A3]=8'h00;
    mem['h52A4]=8'h00; mem['h52A5]=8'h00; mem['h52A6]=8'h00; mem['h52A7]=8'h00;
    mem['h52A8]=8'h00; mem['h52A9]=8'h00; mem['h52AA]=8'h00; mem['h52AB]=8'h00;
    mem['h52AC]=8'h00; mem['h52AD]=8'h00; mem['h52AE]=8'h00; mem['h52AF]=8'h00;
    mem['h52B0]=8'h00; mem['h52B1]=8'h00; mem['h52B2]=8'h00; mem['h52B3]=8'h00;
    mem['h52B4]=8'h00; mem['h52B5]=8'h00; mem['h52B6]=8'h00; mem['h52B7]=8'h00;
    mem['h52B8]=8'h00; mem['h52B9]=8'h00; mem['h52BA]=8'h00; mem['h52BB]=8'h00;
    mem['h52BC]=8'h00; mem['h52BD]=8'h00; mem['h52BE]=8'h00; mem['h52BF]=8'h00;
    mem['h52C0]=8'h00; mem['h52C1]=8'h00; mem['h52C2]=8'h00; mem['h52C3]=8'h00;
    mem['h52C4]=8'h00; mem['h52C5]=8'h00; mem['h52C6]=8'h00; mem['h52C7]=8'h00;
    mem['h52C8]=8'h00; mem['h52C9]=8'h00; mem['h52CA]=8'h00; mem['h52CB]=8'h00;
    mem['h52CC]=8'h00; mem['h52CD]=8'h00; mem['h52CE]=8'h00; mem['h52CF]=8'h00;
    mem['h52D0]=8'h00; mem['h52D1]=8'h00; mem['h52D2]=8'h00; mem['h52D3]=8'h00;
    mem['h52D4]=8'h00; mem['h52D5]=8'h00; mem['h52D6]=8'h00; mem['h52D7]=8'h00;
    mem['h52D8]=8'h00; mem['h52D9]=8'h00; mem['h52DA]=8'h00; mem['h52DB]=8'h00;
    mem['h52DC]=8'h00; mem['h52DD]=8'h00; mem['h52DE]=8'h00; mem['h52DF]=8'h00;
    mem['h52E0]=8'h00; mem['h52E1]=8'h00; mem['h52E2]=8'h00; mem['h52E3]=8'h00;
    mem['h52E4]=8'h00; mem['h52E5]=8'h00; mem['h52E6]=8'h00; mem['h52E7]=8'h00;
    mem['h52E8]=8'h00; mem['h52E9]=8'h00; mem['h52EA]=8'h00; mem['h52EB]=8'h00;
    mem['h52EC]=8'h00; mem['h52ED]=8'h00; mem['h52EE]=8'h00; mem['h52EF]=8'h00;
    mem['h52F0]=8'h00; mem['h52F1]=8'h00; mem['h52F2]=8'h00; mem['h52F3]=8'h00;
    mem['h52F4]=8'h00; mem['h52F5]=8'h00; mem['h52F6]=8'h00; mem['h52F7]=8'h00;
    mem['h52F8]=8'h00; mem['h52F9]=8'h00; mem['h52FA]=8'h00; mem['h52FB]=8'h00;
    mem['h52FC]=8'h00; mem['h52FD]=8'h00; mem['h52FE]=8'h00; mem['h52FF]=8'h00;
    mem['h5300]=8'h00; mem['h5301]=8'h00; mem['h5302]=8'h00; mem['h5303]=8'h00;
    mem['h5304]=8'h00; mem['h5305]=8'h00; mem['h5306]=8'h00; mem['h5307]=8'h00;
    mem['h5308]=8'h00; mem['h5309]=8'h00; mem['h530A]=8'h00; mem['h530B]=8'h00;
    mem['h530C]=8'h00; mem['h530D]=8'h00; mem['h530E]=8'h00; mem['h530F]=8'h00;
    mem['h5310]=8'h00; mem['h5311]=8'h00; mem['h5312]=8'h00; mem['h5313]=8'h00;
    mem['h5314]=8'h00; mem['h5315]=8'h00; mem['h5316]=8'h00; mem['h5317]=8'h00;
    mem['h5318]=8'h00; mem['h5319]=8'h00; mem['h531A]=8'h00; mem['h531B]=8'h00;
    mem['h531C]=8'h00; mem['h531D]=8'h00; mem['h531E]=8'h00; mem['h531F]=8'h00;
    mem['h5320]=8'h00; mem['h5321]=8'h00; mem['h5322]=8'h00; mem['h5323]=8'h00;
    mem['h5324]=8'h00; mem['h5325]=8'h00; mem['h5326]=8'h00; mem['h5327]=8'h00;
    mem['h5328]=8'h00; mem['h5329]=8'h00; mem['h532A]=8'h00; mem['h532B]=8'h00;
    mem['h532C]=8'h00; mem['h532D]=8'h00; mem['h532E]=8'h00; mem['h532F]=8'h00;
    mem['h5330]=8'h00; mem['h5331]=8'h00; mem['h5332]=8'h00; mem['h5333]=8'h00;
    mem['h5334]=8'h00; mem['h5335]=8'h00; mem['h5336]=8'h00; mem['h5337]=8'h00;
    mem['h5338]=8'h00; mem['h5339]=8'h00; mem['h533A]=8'h00; mem['h533B]=8'h00;
    mem['h533C]=8'h00; mem['h533D]=8'h00; mem['h533E]=8'h00; mem['h533F]=8'h00;
    mem['h5340]=8'h00; mem['h5341]=8'h00; mem['h5342]=8'h00; mem['h5343]=8'h00;
    mem['h5344]=8'h00; mem['h5345]=8'h00; mem['h5346]=8'h00; mem['h5347]=8'h00;
    mem['h5348]=8'h00; mem['h5349]=8'h00; mem['h534A]=8'h00; mem['h534B]=8'h00;
    mem['h534C]=8'h00; mem['h534D]=8'h00; mem['h534E]=8'h00; mem['h534F]=8'h00;
    mem['h5350]=8'h00; mem['h5351]=8'h00; mem['h5352]=8'h00; mem['h5353]=8'h00;
    mem['h5354]=8'h00; mem['h5355]=8'h00; mem['h5356]=8'h00; mem['h5357]=8'h00;
    mem['h5358]=8'h00; mem['h5359]=8'h00; mem['h535A]=8'h00; mem['h535B]=8'h00;
    mem['h535C]=8'h00; mem['h535D]=8'h00; mem['h535E]=8'h00; mem['h535F]=8'h00;
    mem['h5360]=8'h00; mem['h5361]=8'h00; mem['h5362]=8'h00; mem['h5363]=8'h00;
    mem['h5364]=8'h00; mem['h5365]=8'h00; mem['h5366]=8'h00; mem['h5367]=8'h00;
    mem['h5368]=8'h00; mem['h5369]=8'h00; mem['h536A]=8'h00; mem['h536B]=8'h00;
    mem['h536C]=8'h00; mem['h536D]=8'h00; mem['h536E]=8'h00; mem['h536F]=8'h00;
    mem['h5370]=8'h00; mem['h5371]=8'h00; mem['h5372]=8'h00; mem['h5373]=8'h00;
    mem['h5374]=8'h00; mem['h5375]=8'h00; mem['h5376]=8'h00; mem['h5377]=8'h00;
    mem['h5378]=8'h00; mem['h5379]=8'h00; mem['h537A]=8'h00; mem['h537B]=8'h00;
    mem['h537C]=8'h00; mem['h537D]=8'h00; mem['h537E]=8'h00; mem['h537F]=8'h00;
    mem['h5380]=8'h00; mem['h5381]=8'h00; mem['h5382]=8'h00; mem['h5383]=8'h00;
    mem['h5384]=8'h00; mem['h5385]=8'h00; mem['h5386]=8'h00; mem['h5387]=8'h00;
    mem['h5388]=8'h00; mem['h5389]=8'h00; mem['h538A]=8'h00; mem['h538B]=8'h00;
    mem['h538C]=8'h00; mem['h538D]=8'h00; mem['h538E]=8'h00; mem['h538F]=8'h00;
    mem['h5390]=8'h00; mem['h5391]=8'h00; mem['h5392]=8'h00; mem['h5393]=8'h00;
    mem['h5394]=8'h00; mem['h5395]=8'h00; mem['h5396]=8'h00; mem['h5397]=8'h00;
    mem['h5398]=8'h00; mem['h5399]=8'h00; mem['h539A]=8'h00; mem['h539B]=8'h00;
    mem['h539C]=8'h00; mem['h539D]=8'h00; mem['h539E]=8'h00; mem['h539F]=8'h00;
    mem['h53A0]=8'h00; mem['h53A1]=8'h00; mem['h53A2]=8'h00; mem['h53A3]=8'h00;
    mem['h53A4]=8'h00; mem['h53A5]=8'h00; mem['h53A6]=8'h00; mem['h53A7]=8'h00;
    mem['h53A8]=8'h00; mem['h53A9]=8'h00; mem['h53AA]=8'h00; mem['h53AB]=8'h00;
    mem['h53AC]=8'h00; mem['h53AD]=8'h00; mem['h53AE]=8'h00; mem['h53AF]=8'h00;
    mem['h53B0]=8'h00; mem['h53B1]=8'h00; mem['h53B2]=8'h00; mem['h53B3]=8'h00;
    mem['h53B4]=8'h00; mem['h53B5]=8'h00; mem['h53B6]=8'h00; mem['h53B7]=8'h00;
    mem['h53B8]=8'h00; mem['h53B9]=8'h00; mem['h53BA]=8'h00; mem['h53BB]=8'h00;
    mem['h53BC]=8'h00; mem['h53BD]=8'h00; mem['h53BE]=8'h00; mem['h53BF]=8'h00;
    mem['h53C0]=8'h00; mem['h53C1]=8'h00; mem['h53C2]=8'h00; mem['h53C3]=8'h00;
    mem['h53C4]=8'h00; mem['h53C5]=8'h00; mem['h53C6]=8'h00; mem['h53C7]=8'h00;
    mem['h53C8]=8'h00; mem['h53C9]=8'h00; mem['h53CA]=8'h00; mem['h53CB]=8'h00;
    mem['h53CC]=8'h00; mem['h53CD]=8'h00; mem['h53CE]=8'h00; mem['h53CF]=8'h00;
    mem['h53D0]=8'h00; mem['h53D1]=8'h00; mem['h53D2]=8'h00; mem['h53D3]=8'h00;
    mem['h53D4]=8'h00; mem['h53D5]=8'h00; mem['h53D6]=8'h00; mem['h53D7]=8'h00;
    mem['h53D8]=8'h00; mem['h53D9]=8'h00; mem['h53DA]=8'h00; mem['h53DB]=8'h00;
    mem['h53DC]=8'h00; mem['h53DD]=8'h00; mem['h53DE]=8'h00; mem['h53DF]=8'h00;
    mem['h53E0]=8'h00; mem['h53E1]=8'h00; mem['h53E2]=8'h00; mem['h53E3]=8'h00;
    mem['h53E4]=8'h00; mem['h53E5]=8'h00; mem['h53E6]=8'h00; mem['h53E7]=8'h00;
    mem['h53E8]=8'h00; mem['h53E9]=8'h00; mem['h53EA]=8'h00; mem['h53EB]=8'h00;
    mem['h53EC]=8'h00; mem['h53ED]=8'h00; mem['h53EE]=8'h00; mem['h53EF]=8'h00;
    mem['h53F0]=8'h00; mem['h53F1]=8'h00; mem['h53F2]=8'h00; mem['h53F3]=8'h00;
    mem['h53F4]=8'h00; mem['h53F5]=8'h00; mem['h53F6]=8'h00; mem['h53F7]=8'h00;
    mem['h53F8]=8'h00; mem['h53F9]=8'h00; mem['h53FA]=8'h00; mem['h53FB]=8'h00;
    mem['h53FC]=8'h00; mem['h53FD]=8'h00; mem['h53FE]=8'h00; mem['h53FF]=8'h00;
    mem['h5400]=8'h00; mem['h5401]=8'h00; mem['h5402]=8'h00; mem['h5403]=8'h00;
    mem['h5404]=8'h00; mem['h5405]=8'h00; mem['h5406]=8'h00; mem['h5407]=8'h00;
    mem['h5408]=8'h00; mem['h5409]=8'h00; mem['h540A]=8'h00; mem['h540B]=8'h00;
    mem['h540C]=8'h00; mem['h540D]=8'h00; mem['h540E]=8'h00; mem['h540F]=8'h00;
    mem['h5410]=8'h00; mem['h5411]=8'h00; mem['h5412]=8'h00; mem['h5413]=8'h00;
    mem['h5414]=8'h00; mem['h5415]=8'h00; mem['h5416]=8'h00; mem['h5417]=8'h00;
    mem['h5418]=8'h00; mem['h5419]=8'h00; mem['h541A]=8'h00; mem['h541B]=8'h00;
    mem['h541C]=8'h00; mem['h541D]=8'h00; mem['h541E]=8'h00; mem['h541F]=8'h00;
    mem['h5420]=8'h00; mem['h5421]=8'h00; mem['h5422]=8'h00; mem['h5423]=8'h00;
    mem['h5424]=8'h00; mem['h5425]=8'h00; mem['h5426]=8'h00; mem['h5427]=8'h00;
    mem['h5428]=8'h00; mem['h5429]=8'h00; mem['h542A]=8'h00; mem['h542B]=8'h00;
    mem['h542C]=8'h00; mem['h542D]=8'h00; mem['h542E]=8'h00; mem['h542F]=8'h00;
    mem['h5430]=8'h00; mem['h5431]=8'h00; mem['h5432]=8'h00; mem['h5433]=8'h00;
    mem['h5434]=8'h00; mem['h5435]=8'h00; mem['h5436]=8'h00; mem['h5437]=8'h00;
    mem['h5438]=8'h00; mem['h5439]=8'h00; mem['h543A]=8'h00; mem['h543B]=8'h00;
    mem['h543C]=8'h00; mem['h543D]=8'h00; mem['h543E]=8'h00; mem['h543F]=8'h00;
    mem['h5440]=8'h00; mem['h5441]=8'h00; mem['h5442]=8'h00; mem['h5443]=8'h00;
    mem['h5444]=8'h00; mem['h5445]=8'h00; mem['h5446]=8'h00; mem['h5447]=8'h00;
    mem['h5448]=8'h00; mem['h5449]=8'h00; mem['h544A]=8'h00; mem['h544B]=8'h00;
    mem['h544C]=8'h00; mem['h544D]=8'h00; mem['h544E]=8'h00; mem['h544F]=8'h00;
    mem['h5450]=8'h00; mem['h5451]=8'h00; mem['h5452]=8'h00; mem['h5453]=8'h00;
    mem['h5454]=8'h00; mem['h5455]=8'h00; mem['h5456]=8'h00; mem['h5457]=8'h00;
    mem['h5458]=8'h00; mem['h5459]=8'h00; mem['h545A]=8'h00; mem['h545B]=8'h00;
    mem['h545C]=8'h00; mem['h545D]=8'h00; mem['h545E]=8'h00; mem['h545F]=8'h00;
    mem['h5460]=8'h00; mem['h5461]=8'h00; mem['h5462]=8'h00; mem['h5463]=8'h00;
    mem['h5464]=8'h00; mem['h5465]=8'h00; mem['h5466]=8'h00; mem['h5467]=8'h00;
    mem['h5468]=8'h00; mem['h5469]=8'h00; mem['h546A]=8'h00; mem['h546B]=8'h00;
    mem['h546C]=8'h00; mem['h546D]=8'h00; mem['h546E]=8'h00; mem['h546F]=8'h00;
    mem['h5470]=8'h00; mem['h5471]=8'h00; mem['h5472]=8'h00; mem['h5473]=8'h00;
    mem['h5474]=8'h00; mem['h5475]=8'h00; mem['h5476]=8'h00; mem['h5477]=8'h00;
    mem['h5478]=8'h00; mem['h5479]=8'h00; mem['h547A]=8'h00; mem['h547B]=8'h00;
    mem['h547C]=8'h00; mem['h547D]=8'h00; mem['h547E]=8'h00; mem['h547F]=8'h00;
    mem['h5480]=8'h00; mem['h5481]=8'h00; mem['h5482]=8'h00; mem['h5483]=8'h00;
    mem['h5484]=8'h00; mem['h5485]=8'h00; mem['h5486]=8'h00; mem['h5487]=8'h00;
    mem['h5488]=8'h00; mem['h5489]=8'h00; mem['h548A]=8'h00; mem['h548B]=8'h00;
    mem['h548C]=8'h00; mem['h548D]=8'h00; mem['h548E]=8'h00; mem['h548F]=8'h00;
    mem['h5490]=8'h00; mem['h5491]=8'h00; mem['h5492]=8'h00; mem['h5493]=8'h00;
    mem['h5494]=8'h00; mem['h5495]=8'h00; mem['h5496]=8'h00; mem['h5497]=8'h00;
    mem['h5498]=8'h00; mem['h5499]=8'h00; mem['h549A]=8'h00; mem['h549B]=8'h00;
    mem['h549C]=8'h00; mem['h549D]=8'h00; mem['h549E]=8'h00; mem['h549F]=8'h00;
    mem['h54A0]=8'h00; mem['h54A1]=8'h00; mem['h54A2]=8'h00; mem['h54A3]=8'h00;
    mem['h54A4]=8'h00; mem['h54A5]=8'h00; mem['h54A6]=8'h00; mem['h54A7]=8'h00;
    mem['h54A8]=8'h00; mem['h54A9]=8'h00; mem['h54AA]=8'h00; mem['h54AB]=8'h00;
    mem['h54AC]=8'h00; mem['h54AD]=8'h00; mem['h54AE]=8'h00; mem['h54AF]=8'h00;
    mem['h54B0]=8'h00; mem['h54B1]=8'h00; mem['h54B2]=8'h00; mem['h54B3]=8'h00;
    mem['h54B4]=8'h00; mem['h54B5]=8'h00; mem['h54B6]=8'h00; mem['h54B7]=8'h00;
    mem['h54B8]=8'h00; mem['h54B9]=8'h00; mem['h54BA]=8'h00; mem['h54BB]=8'h00;
    mem['h54BC]=8'h00; mem['h54BD]=8'h00; mem['h54BE]=8'h00; mem['h54BF]=8'h00;
    mem['h54C0]=8'h00; mem['h54C1]=8'h00; mem['h54C2]=8'h00; mem['h54C3]=8'h00;
    mem['h54C4]=8'h00; mem['h54C5]=8'h00; mem['h54C6]=8'h00; mem['h54C7]=8'h00;
    mem['h54C8]=8'h00; mem['h54C9]=8'h00; mem['h54CA]=8'h00; mem['h54CB]=8'h00;
    mem['h54CC]=8'h00; mem['h54CD]=8'h00; mem['h54CE]=8'h00; mem['h54CF]=8'h00;
    mem['h54D0]=8'h00; mem['h54D1]=8'h00; mem['h54D2]=8'h00; mem['h54D3]=8'h00;
    mem['h54D4]=8'h00; mem['h54D5]=8'h00; mem['h54D6]=8'h00; mem['h54D7]=8'h00;
    mem['h54D8]=8'h00; mem['h54D9]=8'h00; mem['h54DA]=8'h00; mem['h54DB]=8'h00;
    mem['h54DC]=8'h00; mem['h54DD]=8'h00; mem['h54DE]=8'h00; mem['h54DF]=8'h00;
    mem['h54E0]=8'h00; mem['h54E1]=8'h00; mem['h54E2]=8'h00; mem['h54E3]=8'h00;
    mem['h54E4]=8'h00; mem['h54E5]=8'h00; mem['h54E6]=8'h00; mem['h54E7]=8'h00;
    mem['h54E8]=8'h00; mem['h54E9]=8'h00; mem['h54EA]=8'h00; mem['h54EB]=8'h00;
    mem['h54EC]=8'h00; mem['h54ED]=8'h00; mem['h54EE]=8'h00; mem['h54EF]=8'h00;
    mem['h54F0]=8'h00; mem['h54F1]=8'h00; mem['h54F2]=8'h00; mem['h54F3]=8'h00;
    mem['h54F4]=8'h00; mem['h54F5]=8'h00; mem['h54F6]=8'h00; mem['h54F7]=8'h00;
    mem['h54F8]=8'h00; mem['h54F9]=8'h00; mem['h54FA]=8'h00; mem['h54FB]=8'h00;
    mem['h54FC]=8'h00; mem['h54FD]=8'h00; mem['h54FE]=8'h00; mem['h54FF]=8'h00;
    mem['h5500]=8'h00; mem['h5501]=8'h00; mem['h5502]=8'h00; mem['h5503]=8'h00;
    mem['h5504]=8'h00; mem['h5505]=8'h00; mem['h5506]=8'h00; mem['h5507]=8'h00;
    mem['h5508]=8'h00; mem['h5509]=8'h00; mem['h550A]=8'h00; mem['h550B]=8'h00;
    mem['h550C]=8'h00; mem['h550D]=8'h00; mem['h550E]=8'h00; mem['h550F]=8'h00;
    mem['h5510]=8'h00; mem['h5511]=8'h00; mem['h5512]=8'h00; mem['h5513]=8'h00;
    mem['h5514]=8'h00; mem['h5515]=8'h00; mem['h5516]=8'h00; mem['h5517]=8'h00;
    mem['h5518]=8'h00; mem['h5519]=8'h00; mem['h551A]=8'h00; mem['h551B]=8'h00;
    mem['h551C]=8'h00; mem['h551D]=8'h00; mem['h551E]=8'h00; mem['h551F]=8'h00;
    mem['h5520]=8'h00; mem['h5521]=8'h00; mem['h5522]=8'h00; mem['h5523]=8'h00;
    mem['h5524]=8'h00; mem['h5525]=8'h00; mem['h5526]=8'h00; mem['h5527]=8'h00;
    mem['h5528]=8'h00; mem['h5529]=8'h00; mem['h552A]=8'h00; mem['h552B]=8'h00;
    mem['h552C]=8'h00; mem['h552D]=8'h00; mem['h552E]=8'h00; mem['h552F]=8'h00;
    mem['h5530]=8'h00; mem['h5531]=8'h00; mem['h5532]=8'h00; mem['h5533]=8'h00;
    mem['h5534]=8'h00; mem['h5535]=8'h00; mem['h5536]=8'h00; mem['h5537]=8'h00;
    mem['h5538]=8'h00; mem['h5539]=8'h00; mem['h553A]=8'h00; mem['h553B]=8'h00;
    mem['h553C]=8'h00; mem['h553D]=8'h00; mem['h553E]=8'h00; mem['h553F]=8'h00;
    mem['h5540]=8'h00; mem['h5541]=8'h00; mem['h5542]=8'h00; mem['h5543]=8'h00;
    mem['h5544]=8'h00; mem['h5545]=8'h00; mem['h5546]=8'h00; mem['h5547]=8'h00;
    mem['h5548]=8'h00; mem['h5549]=8'h00; mem['h554A]=8'h00; mem['h554B]=8'h00;
    mem['h554C]=8'h00; mem['h554D]=8'h00; mem['h554E]=8'h00; mem['h554F]=8'h00;
    mem['h5550]=8'h00; mem['h5551]=8'h00; mem['h5552]=8'h00; mem['h5553]=8'h00;
    mem['h5554]=8'h00; mem['h5555]=8'h00; mem['h5556]=8'h00; mem['h5557]=8'h00;
    mem['h5558]=8'h00; mem['h5559]=8'h00; mem['h555A]=8'h00; mem['h555B]=8'h00;
    mem['h555C]=8'h00; mem['h555D]=8'h00; mem['h555E]=8'h00; mem['h555F]=8'h00;
    mem['h5560]=8'h00; mem['h5561]=8'h00; mem['h5562]=8'h00; mem['h5563]=8'h00;
    mem['h5564]=8'h00; mem['h5565]=8'h00; mem['h5566]=8'h00; mem['h5567]=8'h00;
    mem['h5568]=8'h00; mem['h5569]=8'h00; mem['h556A]=8'h00; mem['h556B]=8'h00;
    mem['h556C]=8'h00; mem['h556D]=8'h00; mem['h556E]=8'h00; mem['h556F]=8'h00;
    mem['h5570]=8'h00; mem['h5571]=8'h00; mem['h5572]=8'h00; mem['h5573]=8'h00;
    mem['h5574]=8'h00; mem['h5575]=8'h00; mem['h5576]=8'h00; mem['h5577]=8'h00;
    mem['h5578]=8'h00; mem['h5579]=8'h00; mem['h557A]=8'h00; mem['h557B]=8'h00;
    mem['h557C]=8'h00; mem['h557D]=8'h00; mem['h557E]=8'h00; mem['h557F]=8'h00;
    mem['h5580]=8'h00; mem['h5581]=8'h00; mem['h5582]=8'h00; mem['h5583]=8'h00;
    mem['h5584]=8'h00; mem['h5585]=8'h00; mem['h5586]=8'h00; mem['h5587]=8'h00;
    mem['h5588]=8'h00; mem['h5589]=8'h00; mem['h558A]=8'h00; mem['h558B]=8'h00;
    mem['h558C]=8'h00; mem['h558D]=8'h00; mem['h558E]=8'h00; mem['h558F]=8'h00;
    mem['h5590]=8'h00; mem['h5591]=8'h00; mem['h5592]=8'h00; mem['h5593]=8'h00;
    mem['h5594]=8'h00; mem['h5595]=8'h00; mem['h5596]=8'h00; mem['h5597]=8'h00;
    mem['h5598]=8'h00; mem['h5599]=8'h00; mem['h559A]=8'h00; mem['h559B]=8'h00;
    mem['h559C]=8'h00; mem['h559D]=8'h00; mem['h559E]=8'h00; mem['h559F]=8'h00;
    mem['h55A0]=8'h00; mem['h55A1]=8'h00; mem['h55A2]=8'h00; mem['h55A3]=8'h00;
    mem['h55A4]=8'h00; mem['h55A5]=8'h00; mem['h55A6]=8'h00; mem['h55A7]=8'h00;
    mem['h55A8]=8'h00; mem['h55A9]=8'h00; mem['h55AA]=8'h00; mem['h55AB]=8'h00;
    mem['h55AC]=8'h00; mem['h55AD]=8'h00; mem['h55AE]=8'h00; mem['h55AF]=8'h00;
    mem['h55B0]=8'h00; mem['h55B1]=8'h00; mem['h55B2]=8'h00; mem['h55B3]=8'h00;
    mem['h55B4]=8'h00; mem['h55B5]=8'h00; mem['h55B6]=8'h00; mem['h55B7]=8'h00;
    mem['h55B8]=8'h00; mem['h55B9]=8'h00; mem['h55BA]=8'h00; mem['h55BB]=8'h00;
    mem['h55BC]=8'h00; mem['h55BD]=8'h00; mem['h55BE]=8'h00; mem['h55BF]=8'h00;
    mem['h55C0]=8'h00; mem['h55C1]=8'h00; mem['h55C2]=8'h00; mem['h55C3]=8'h00;
    mem['h55C4]=8'h00; mem['h55C5]=8'h00; mem['h55C6]=8'h00; mem['h55C7]=8'h00;
    mem['h55C8]=8'h00; mem['h55C9]=8'h00; mem['h55CA]=8'h00; mem['h55CB]=8'h00;
    mem['h55CC]=8'h00; mem['h55CD]=8'h00; mem['h55CE]=8'h00; mem['h55CF]=8'h00;
    mem['h55D0]=8'h00; mem['h55D1]=8'h00; mem['h55D2]=8'h00; mem['h55D3]=8'h00;
    mem['h55D4]=8'h00; mem['h55D5]=8'h00; mem['h55D6]=8'h00; mem['h55D7]=8'h00;
    mem['h55D8]=8'h00; mem['h55D9]=8'h00; mem['h55DA]=8'h00; mem['h55DB]=8'h00;
    mem['h55DC]=8'h00; mem['h55DD]=8'h00; mem['h55DE]=8'h00; mem['h55DF]=8'h00;
    mem['h55E0]=8'h00; mem['h55E1]=8'h00; mem['h55E2]=8'h00; mem['h55E3]=8'h00;
    mem['h55E4]=8'h00; mem['h55E5]=8'h00; mem['h55E6]=8'h00; mem['h55E7]=8'h00;
    mem['h55E8]=8'h00; mem['h55E9]=8'h00; mem['h55EA]=8'h00; mem['h55EB]=8'h00;
    mem['h55EC]=8'h00; mem['h55ED]=8'h00; mem['h55EE]=8'h00; mem['h55EF]=8'h00;
    mem['h55F0]=8'h00; mem['h55F1]=8'h00; mem['h55F2]=8'h00; mem['h55F3]=8'h00;
    mem['h55F4]=8'h00; mem['h55F5]=8'h00; mem['h55F6]=8'h00; mem['h55F7]=8'h00;
    mem['h55F8]=8'h00; mem['h55F9]=8'h00; mem['h55FA]=8'h00; mem['h55FB]=8'h00;
    mem['h55FC]=8'h00; mem['h55FD]=8'h00; mem['h55FE]=8'h00; mem['h55FF]=8'h00;
    mem['h5600]=8'h00; mem['h5601]=8'h00; mem['h5602]=8'h00; mem['h5603]=8'h00;
    mem['h5604]=8'h00; mem['h5605]=8'h00; mem['h5606]=8'h00; mem['h5607]=8'h00;
    mem['h5608]=8'h00; mem['h5609]=8'h00; mem['h560A]=8'h00; mem['h560B]=8'h00;
    mem['h560C]=8'h00; mem['h560D]=8'h00; mem['h560E]=8'h00; mem['h560F]=8'h00;
    mem['h5610]=8'h00; mem['h5611]=8'h00; mem['h5612]=8'h00; mem['h5613]=8'h00;
    mem['h5614]=8'h00; mem['h5615]=8'h00; mem['h5616]=8'h00; mem['h5617]=8'h00;
    mem['h5618]=8'h00; mem['h5619]=8'h00; mem['h561A]=8'h00; mem['h561B]=8'h00;
    mem['h561C]=8'h00; mem['h561D]=8'h00; mem['h561E]=8'h00; mem['h561F]=8'h00;
    mem['h5620]=8'h00; mem['h5621]=8'h00; mem['h5622]=8'h00; mem['h5623]=8'h00;
    mem['h5624]=8'h00; mem['h5625]=8'h00; mem['h5626]=8'h00; mem['h5627]=8'h00;
    mem['h5628]=8'h00; mem['h5629]=8'h00; mem['h562A]=8'h00; mem['h562B]=8'h00;
    mem['h562C]=8'h00; mem['h562D]=8'h00; mem['h562E]=8'h00; mem['h562F]=8'h00;
    mem['h5630]=8'h00; mem['h5631]=8'h00; mem['h5632]=8'h00; mem['h5633]=8'h00;
    mem['h5634]=8'h00; mem['h5635]=8'h00; mem['h5636]=8'h00; mem['h5637]=8'h00;
    mem['h5638]=8'h00; mem['h5639]=8'h00; mem['h563A]=8'h00; mem['h563B]=8'h00;
    mem['h563C]=8'h00; mem['h563D]=8'h00; mem['h563E]=8'h00; mem['h563F]=8'h00;
    mem['h5640]=8'h00; mem['h5641]=8'h00; mem['h5642]=8'h00; mem['h5643]=8'h00;
    mem['h5644]=8'h00; mem['h5645]=8'h00; mem['h5646]=8'h00; mem['h5647]=8'h00;
    mem['h5648]=8'h00; mem['h5649]=8'h00; mem['h564A]=8'h00; mem['h564B]=8'h00;
    mem['h564C]=8'h00; mem['h564D]=8'h00; mem['h564E]=8'h00; mem['h564F]=8'h00;
    mem['h5650]=8'h00; mem['h5651]=8'h00; mem['h5652]=8'h00; mem['h5653]=8'h00;
    mem['h5654]=8'h00; mem['h5655]=8'h00; mem['h5656]=8'h00; mem['h5657]=8'h00;
    mem['h5658]=8'h00; mem['h5659]=8'h00; mem['h565A]=8'h00; mem['h565B]=8'h00;
    mem['h565C]=8'h00; mem['h565D]=8'h00; mem['h565E]=8'h00; mem['h565F]=8'h00;
    mem['h5660]=8'h00; mem['h5661]=8'h00; mem['h5662]=8'h00; mem['h5663]=8'h00;
    mem['h5664]=8'h00; mem['h5665]=8'h00; mem['h5666]=8'h00; mem['h5667]=8'h00;
    mem['h5668]=8'h00; mem['h5669]=8'h00; mem['h566A]=8'h00; mem['h566B]=8'h00;
    mem['h566C]=8'h00; mem['h566D]=8'h00; mem['h566E]=8'h00; mem['h566F]=8'h00;
    mem['h5670]=8'h00; mem['h5671]=8'h00; mem['h5672]=8'h00; mem['h5673]=8'h00;
    mem['h5674]=8'h00; mem['h5675]=8'h00; mem['h5676]=8'h00; mem['h5677]=8'h00;
    mem['h5678]=8'h00; mem['h5679]=8'h00; mem['h567A]=8'h00; mem['h567B]=8'h00;
    mem['h567C]=8'h00; mem['h567D]=8'h00; mem['h567E]=8'h00; mem['h567F]=8'h00;
    mem['h5680]=8'h00; mem['h5681]=8'h00; mem['h5682]=8'h00; mem['h5683]=8'h00;
    mem['h5684]=8'h00; mem['h5685]=8'h00; mem['h5686]=8'h00; mem['h5687]=8'h00;
    mem['h5688]=8'h00; mem['h5689]=8'h00; mem['h568A]=8'h00; mem['h568B]=8'h00;
    mem['h568C]=8'h00; mem['h568D]=8'h00; mem['h568E]=8'h00; mem['h568F]=8'h00;
    mem['h5690]=8'h00; mem['h5691]=8'h00; mem['h5692]=8'h00; mem['h5693]=8'h00;
    mem['h5694]=8'h00; mem['h5695]=8'h00; mem['h5696]=8'h00; mem['h5697]=8'h00;
    mem['h5698]=8'h00; mem['h5699]=8'h00; mem['h569A]=8'h00; mem['h569B]=8'h00;
    mem['h569C]=8'h00; mem['h569D]=8'h00; mem['h569E]=8'h00; mem['h569F]=8'h00;
    mem['h56A0]=8'h00; mem['h56A1]=8'h00; mem['h56A2]=8'h00; mem['h56A3]=8'h00;
    mem['h56A4]=8'h00; mem['h56A5]=8'h00; mem['h56A6]=8'h00; mem['h56A7]=8'h00;
    mem['h56A8]=8'h00; mem['h56A9]=8'h00; mem['h56AA]=8'h00; mem['h56AB]=8'h00;
    mem['h56AC]=8'h00; mem['h56AD]=8'h00; mem['h56AE]=8'h00; mem['h56AF]=8'h00;
    mem['h56B0]=8'h00; mem['h56B1]=8'h00; mem['h56B2]=8'h00; mem['h56B3]=8'h00;
    mem['h56B4]=8'h00; mem['h56B5]=8'h00; mem['h56B6]=8'h00; mem['h56B7]=8'h00;
    mem['h56B8]=8'h00; mem['h56B9]=8'h00; mem['h56BA]=8'h00; mem['h56BB]=8'h00;
    mem['h56BC]=8'h00; mem['h56BD]=8'h00; mem['h56BE]=8'h00; mem['h56BF]=8'h00;
    mem['h56C0]=8'h00; mem['h56C1]=8'h00; mem['h56C2]=8'h00; mem['h56C3]=8'h00;
    mem['h56C4]=8'h00; mem['h56C5]=8'h00; mem['h56C6]=8'h00; mem['h56C7]=8'h00;
    mem['h56C8]=8'h00; mem['h56C9]=8'h00; mem['h56CA]=8'h00; mem['h56CB]=8'h00;
    mem['h56CC]=8'h00; mem['h56CD]=8'h00; mem['h56CE]=8'h00; mem['h56CF]=8'h00;
    mem['h56D0]=8'h00; mem['h56D1]=8'h00; mem['h56D2]=8'h00; mem['h56D3]=8'h00;
    mem['h56D4]=8'h00; mem['h56D5]=8'h00; mem['h56D6]=8'h00; mem['h56D7]=8'h00;
    mem['h56D8]=8'h00; mem['h56D9]=8'h00; mem['h56DA]=8'h00; mem['h56DB]=8'h00;
    mem['h56DC]=8'h00; mem['h56DD]=8'h00; mem['h56DE]=8'h00; mem['h56DF]=8'h00;
    mem['h56E0]=8'h00; mem['h56E1]=8'h00; mem['h56E2]=8'h00; mem['h56E3]=8'h00;
    mem['h56E4]=8'h00; mem['h56E5]=8'h00; mem['h56E6]=8'h00; mem['h56E7]=8'h00;
    mem['h56E8]=8'h00; mem['h56E9]=8'h00; mem['h56EA]=8'h00; mem['h56EB]=8'h00;
    mem['h56EC]=8'h00; mem['h56ED]=8'h00; mem['h56EE]=8'h00; mem['h56EF]=8'h00;
    mem['h56F0]=8'h00; mem['h56F1]=8'h00; mem['h56F2]=8'h00; mem['h56F3]=8'h00;
    mem['h56F4]=8'h00; mem['h56F5]=8'h00; mem['h56F6]=8'h00; mem['h56F7]=8'h00;
    mem['h56F8]=8'h00; mem['h56F9]=8'h00; mem['h56FA]=8'h00; mem['h56FB]=8'h00;
    mem['h56FC]=8'h00; mem['h56FD]=8'h00; mem['h56FE]=8'h00; mem['h56FF]=8'h00;
    mem['h5700]=8'h00; mem['h5701]=8'h00; mem['h5702]=8'h00; mem['h5703]=8'h00;
    mem['h5704]=8'h00; mem['h5705]=8'h00; mem['h5706]=8'h00; mem['h5707]=8'h00;
    mem['h5708]=8'h00; mem['h5709]=8'h00; mem['h570A]=8'h00; mem['h570B]=8'h00;
    mem['h570C]=8'h00; mem['h570D]=8'h00; mem['h570E]=8'h00; mem['h570F]=8'h00;
    mem['h5710]=8'h00; mem['h5711]=8'h00; mem['h5712]=8'h00; mem['h5713]=8'h00;
    mem['h5714]=8'h00; mem['h5715]=8'h00; mem['h5716]=8'h00; mem['h5717]=8'h00;
    mem['h5718]=8'h00; mem['h5719]=8'h00; mem['h571A]=8'h00; mem['h571B]=8'h00;
    mem['h571C]=8'h00; mem['h571D]=8'h00; mem['h571E]=8'h00; mem['h571F]=8'h00;
    mem['h5720]=8'h00; mem['h5721]=8'h00; mem['h5722]=8'h00; mem['h5723]=8'h00;
    mem['h5724]=8'h00; mem['h5725]=8'h00; mem['h5726]=8'h00; mem['h5727]=8'h00;
    mem['h5728]=8'h00; mem['h5729]=8'h00; mem['h572A]=8'h00; mem['h572B]=8'h00;
    mem['h572C]=8'h00; mem['h572D]=8'h00; mem['h572E]=8'h00; mem['h572F]=8'h00;
    mem['h5730]=8'h00; mem['h5731]=8'h00; mem['h5732]=8'h00; mem['h5733]=8'h00;
    mem['h5734]=8'h00; mem['h5735]=8'h00; mem['h5736]=8'h00; mem['h5737]=8'h00;
    mem['h5738]=8'h00; mem['h5739]=8'h00; mem['h573A]=8'h00; mem['h573B]=8'h00;
    mem['h573C]=8'h00; mem['h573D]=8'h00; mem['h573E]=8'h00; mem['h573F]=8'h00;
    mem['h5740]=8'h00; mem['h5741]=8'h00; mem['h5742]=8'h00; mem['h5743]=8'h00;
    mem['h5744]=8'h00; mem['h5745]=8'h00; mem['h5746]=8'h00; mem['h5747]=8'h00;
    mem['h5748]=8'h00; mem['h5749]=8'h00; mem['h574A]=8'h00; mem['h574B]=8'h00;
    mem['h574C]=8'h00; mem['h574D]=8'h00; mem['h574E]=8'h00; mem['h574F]=8'h00;
    mem['h5750]=8'h00; mem['h5751]=8'h00; mem['h5752]=8'h00; mem['h5753]=8'h00;
    mem['h5754]=8'h00; mem['h5755]=8'h00; mem['h5756]=8'h00; mem['h5757]=8'h00;
    mem['h5758]=8'h00; mem['h5759]=8'h00; mem['h575A]=8'h00; mem['h575B]=8'h00;
    mem['h575C]=8'h00; mem['h575D]=8'h00; mem['h575E]=8'h00; mem['h575F]=8'h00;
    mem['h5760]=8'h00; mem['h5761]=8'h00; mem['h5762]=8'h00; mem['h5763]=8'h00;
    mem['h5764]=8'h00; mem['h5765]=8'h00; mem['h5766]=8'h00; mem['h5767]=8'h00;
    mem['h5768]=8'h00; mem['h5769]=8'h00; mem['h576A]=8'h00; mem['h576B]=8'h00;
    mem['h576C]=8'h00; mem['h576D]=8'h00; mem['h576E]=8'h00; mem['h576F]=8'h00;
    mem['h5770]=8'h00; mem['h5771]=8'h00; mem['h5772]=8'h00; mem['h5773]=8'h00;
    mem['h5774]=8'h00; mem['h5775]=8'h00; mem['h5776]=8'h00; mem['h5777]=8'h00;
    mem['h5778]=8'h00; mem['h5779]=8'h00; mem['h577A]=8'h00; mem['h577B]=8'h00;
    mem['h577C]=8'h00; mem['h577D]=8'h00; mem['h577E]=8'h00; mem['h577F]=8'h00;
    mem['h5780]=8'h00; mem['h5781]=8'h00; mem['h5782]=8'h00; mem['h5783]=8'h00;
    mem['h5784]=8'h00; mem['h5785]=8'h00; mem['h5786]=8'h00; mem['h5787]=8'h00;
    mem['h5788]=8'h00; mem['h5789]=8'h00; mem['h578A]=8'h00; mem['h578B]=8'h00;
    mem['h578C]=8'h00; mem['h578D]=8'h00; mem['h578E]=8'h00; mem['h578F]=8'h00;
    mem['h5790]=8'h00; mem['h5791]=8'h00; mem['h5792]=8'h00; mem['h5793]=8'h00;
    mem['h5794]=8'h00; mem['h5795]=8'h00; mem['h5796]=8'h00; mem['h5797]=8'h00;
    mem['h5798]=8'h00; mem['h5799]=8'h00; mem['h579A]=8'h00; mem['h579B]=8'h00;
    mem['h579C]=8'h00; mem['h579D]=8'h00; mem['h579E]=8'h00; mem['h579F]=8'h00;
    mem['h57A0]=8'h00; mem['h57A1]=8'h00; mem['h57A2]=8'h00; mem['h57A3]=8'h00;
    mem['h57A4]=8'h00; mem['h57A5]=8'h00; mem['h57A6]=8'h00; mem['h57A7]=8'h00;
    mem['h57A8]=8'h00; mem['h57A9]=8'h00; mem['h57AA]=8'h00; mem['h57AB]=8'h00;
    mem['h57AC]=8'h00; mem['h57AD]=8'h00; mem['h57AE]=8'h00; mem['h57AF]=8'h00;
    mem['h57B0]=8'h00; mem['h57B1]=8'h00; mem['h57B2]=8'h00; mem['h57B3]=8'h00;
    mem['h57B4]=8'h00; mem['h57B5]=8'h00; mem['h57B6]=8'h00; mem['h57B7]=8'h00;
    mem['h57B8]=8'h00; mem['h57B9]=8'h00; mem['h57BA]=8'h00; mem['h57BB]=8'h00;
    mem['h57BC]=8'h00; mem['h57BD]=8'h00; mem['h57BE]=8'h00; mem['h57BF]=8'h00;
    mem['h57C0]=8'h00; mem['h57C1]=8'h00; mem['h57C2]=8'h00; mem['h57C3]=8'h00;
    mem['h57C4]=8'h00; mem['h57C5]=8'h00; mem['h57C6]=8'h00; mem['h57C7]=8'h00;
    mem['h57C8]=8'h00; mem['h57C9]=8'h00; mem['h57CA]=8'h00; mem['h57CB]=8'h00;
    mem['h57CC]=8'h00; mem['h57CD]=8'h00; mem['h57CE]=8'h00; mem['h57CF]=8'h00;
    mem['h57D0]=8'h00; mem['h57D1]=8'h00; mem['h57D2]=8'h00; mem['h57D3]=8'h00;
    mem['h57D4]=8'h00; mem['h57D5]=8'h00; mem['h57D6]=8'h00; mem['h57D7]=8'h00;
    mem['h57D8]=8'h00; mem['h57D9]=8'h00; mem['h57DA]=8'h00; mem['h57DB]=8'h00;
    mem['h57DC]=8'h00; mem['h57DD]=8'h00; mem['h57DE]=8'h00; mem['h57DF]=8'h00;
    mem['h57E0]=8'h00; mem['h57E1]=8'h00; mem['h57E2]=8'h00; mem['h57E3]=8'h00;
    mem['h57E4]=8'h00; mem['h57E5]=8'h00; mem['h57E6]=8'h00; mem['h57E7]=8'h00;
    mem['h57E8]=8'h00; mem['h57E9]=8'h00; mem['h57EA]=8'h00; mem['h57EB]=8'h00;
    mem['h57EC]=8'h00; mem['h57ED]=8'h00; mem['h57EE]=8'h00; mem['h57EF]=8'h00;
    mem['h57F0]=8'h00; mem['h57F1]=8'h00; mem['h57F2]=8'h00; mem['h57F3]=8'h00;
    mem['h57F4]=8'h00; mem['h57F5]=8'h00; mem['h57F6]=8'h00; mem['h57F7]=8'h00;
    mem['h57F8]=8'h00; mem['h57F9]=8'h00; mem['h57FA]=8'h00; mem['h57FB]=8'h00;
    mem['h57FC]=8'h00; mem['h57FD]=8'h00; mem['h57FE]=8'h00; mem['h57FF]=8'h00;
    mem['h5800]=8'h00; mem['h5801]=8'h00; mem['h5802]=8'h00; mem['h5803]=8'h00;
    mem['h5804]=8'h00; mem['h5805]=8'h00; mem['h5806]=8'h00; mem['h5807]=8'h00;
    mem['h5808]=8'h00; mem['h5809]=8'h00; mem['h580A]=8'h00; mem['h580B]=8'h00;
    mem['h580C]=8'h00; mem['h580D]=8'h00; mem['h580E]=8'h00; mem['h580F]=8'h00;
    mem['h5810]=8'h00; mem['h5811]=8'h00; mem['h5812]=8'h00; mem['h5813]=8'h00;
    mem['h5814]=8'h00; mem['h5815]=8'h00; mem['h5816]=8'h00; mem['h5817]=8'h00;
    mem['h5818]=8'h00; mem['h5819]=8'h00; mem['h581A]=8'h00; mem['h581B]=8'h00;
    mem['h581C]=8'h00; mem['h581D]=8'h00; mem['h581E]=8'h00; mem['h581F]=8'h00;
    mem['h5820]=8'h00; mem['h5821]=8'h00; mem['h5822]=8'h00; mem['h5823]=8'h00;
    mem['h5824]=8'h00; mem['h5825]=8'h00; mem['h5826]=8'h00; mem['h5827]=8'h00;
    mem['h5828]=8'h00; mem['h5829]=8'h00; mem['h582A]=8'h00; mem['h582B]=8'h00;
    mem['h582C]=8'h00; mem['h582D]=8'h00; mem['h582E]=8'h00; mem['h582F]=8'h00;
    mem['h5830]=8'h00; mem['h5831]=8'h00; mem['h5832]=8'h00; mem['h5833]=8'h00;
    mem['h5834]=8'h00; mem['h5835]=8'h00; mem['h5836]=8'h00; mem['h5837]=8'h00;
    mem['h5838]=8'h00; mem['h5839]=8'h00; mem['h583A]=8'h00; mem['h583B]=8'h00;
    mem['h583C]=8'h00; mem['h583D]=8'h00; mem['h583E]=8'h00; mem['h583F]=8'h00;
    mem['h5840]=8'h00; mem['h5841]=8'h00; mem['h5842]=8'h00; mem['h5843]=8'h00;
    mem['h5844]=8'h00; mem['h5845]=8'h00; mem['h5846]=8'h00; mem['h5847]=8'h00;
    mem['h5848]=8'h00; mem['h5849]=8'h00; mem['h584A]=8'h00; mem['h584B]=8'h00;
    mem['h584C]=8'h00; mem['h584D]=8'h00; mem['h584E]=8'h00; mem['h584F]=8'h00;
    mem['h5850]=8'h00; mem['h5851]=8'h00; mem['h5852]=8'h00; mem['h5853]=8'h00;
    mem['h5854]=8'h00; mem['h5855]=8'h00; mem['h5856]=8'h00; mem['h5857]=8'h00;
    mem['h5858]=8'h00; mem['h5859]=8'h00; mem['h585A]=8'h00; mem['h585B]=8'h00;
    mem['h585C]=8'h00; mem['h585D]=8'h00; mem['h585E]=8'h00; mem['h585F]=8'h00;
    mem['h5860]=8'h00; mem['h5861]=8'h00; mem['h5862]=8'h00; mem['h5863]=8'h00;
    mem['h5864]=8'h00; mem['h5865]=8'h00; mem['h5866]=8'h00; mem['h5867]=8'h00;
    mem['h5868]=8'h00; mem['h5869]=8'h00; mem['h586A]=8'h00; mem['h586B]=8'h00;
    mem['h586C]=8'h00; mem['h586D]=8'h00; mem['h586E]=8'h00; mem['h586F]=8'h00;
    mem['h5870]=8'h00; mem['h5871]=8'h00; mem['h5872]=8'h00; mem['h5873]=8'h00;
    mem['h5874]=8'h00; mem['h5875]=8'h00; mem['h5876]=8'h00; mem['h5877]=8'h00;
    mem['h5878]=8'h00; mem['h5879]=8'h00; mem['h587A]=8'h00; mem['h587B]=8'h00;
    mem['h587C]=8'h00; mem['h587D]=8'h00; mem['h587E]=8'h00; mem['h587F]=8'h00;
    mem['h5880]=8'h00; mem['h5881]=8'h00; mem['h5882]=8'h00; mem['h5883]=8'h00;
    mem['h5884]=8'h00; mem['h5885]=8'h00; mem['h5886]=8'h00; mem['h5887]=8'h00;
    mem['h5888]=8'h00; mem['h5889]=8'h00; mem['h588A]=8'h00; mem['h588B]=8'h00;
    mem['h588C]=8'h00; mem['h588D]=8'h00; mem['h588E]=8'h00; mem['h588F]=8'h00;
    mem['h5890]=8'h00; mem['h5891]=8'h00; mem['h5892]=8'h00; mem['h5893]=8'h00;
    mem['h5894]=8'h00; mem['h5895]=8'h00; mem['h5896]=8'h00; mem['h5897]=8'h00;
    mem['h5898]=8'h00; mem['h5899]=8'h00; mem['h589A]=8'h00; mem['h589B]=8'h00;
    mem['h589C]=8'h00; mem['h589D]=8'h00; mem['h589E]=8'h00; mem['h589F]=8'h00;
    mem['h58A0]=8'h00; mem['h58A1]=8'h00; mem['h58A2]=8'h00; mem['h58A3]=8'h00;
    mem['h58A4]=8'h00; mem['h58A5]=8'h00; mem['h58A6]=8'h00; mem['h58A7]=8'h00;
    mem['h58A8]=8'h00; mem['h58A9]=8'h00; mem['h58AA]=8'h00; mem['h58AB]=8'h00;
    mem['h58AC]=8'h00; mem['h58AD]=8'h00; mem['h58AE]=8'h00; mem['h58AF]=8'h00;
    mem['h58B0]=8'h00; mem['h58B1]=8'h00; mem['h58B2]=8'h00; mem['h58B3]=8'h00;
    mem['h58B4]=8'h00; mem['h58B5]=8'h00; mem['h58B6]=8'h00; mem['h58B7]=8'h00;
    mem['h58B8]=8'h00; mem['h58B9]=8'h00; mem['h58BA]=8'h00; mem['h58BB]=8'h00;
    mem['h58BC]=8'h00; mem['h58BD]=8'h00; mem['h58BE]=8'h00; mem['h58BF]=8'h00;
    mem['h58C0]=8'h00; mem['h58C1]=8'h00; mem['h58C2]=8'h00; mem['h58C3]=8'h00;
    mem['h58C4]=8'h00; mem['h58C5]=8'h00; mem['h58C6]=8'h00; mem['h58C7]=8'h00;
    mem['h58C8]=8'h00; mem['h58C9]=8'h00; mem['h58CA]=8'h00; mem['h58CB]=8'h00;
    mem['h58CC]=8'h00; mem['h58CD]=8'h00; mem['h58CE]=8'h00; mem['h58CF]=8'h00;
    mem['h58D0]=8'h00; mem['h58D1]=8'h00; mem['h58D2]=8'h00; mem['h58D3]=8'h00;
    mem['h58D4]=8'h00; mem['h58D5]=8'h00; mem['h58D6]=8'h00; mem['h58D7]=8'h00;
    mem['h58D8]=8'h00; mem['h58D9]=8'h00; mem['h58DA]=8'h00; mem['h58DB]=8'h00;
    mem['h58DC]=8'h00; mem['h58DD]=8'h00; mem['h58DE]=8'h00; mem['h58DF]=8'h00;
    mem['h58E0]=8'h00; mem['h58E1]=8'h00; mem['h58E2]=8'h00; mem['h58E3]=8'h00;
    mem['h58E4]=8'h00; mem['h58E5]=8'h00; mem['h58E6]=8'h00; mem['h58E7]=8'h00;
    mem['h58E8]=8'h00; mem['h58E9]=8'h00; mem['h58EA]=8'h00; mem['h58EB]=8'h00;
    mem['h58EC]=8'h00; mem['h58ED]=8'h00; mem['h58EE]=8'h00; mem['h58EF]=8'h00;
    mem['h58F0]=8'h00; mem['h58F1]=8'h00; mem['h58F2]=8'h00; mem['h58F3]=8'h00;
    mem['h58F4]=8'h00; mem['h58F5]=8'h00; mem['h58F6]=8'h00; mem['h58F7]=8'h00;
    mem['h58F8]=8'h00; mem['h58F9]=8'h00; mem['h58FA]=8'h00; mem['h58FB]=8'h00;
    mem['h58FC]=8'h00; mem['h58FD]=8'h00; mem['h58FE]=8'h00; mem['h58FF]=8'h00;
    mem['h5900]=8'h00; mem['h5901]=8'h00; mem['h5902]=8'h00; mem['h5903]=8'h00;
    mem['h5904]=8'h00; mem['h5905]=8'h00; mem['h5906]=8'h00; mem['h5907]=8'h00;
    mem['h5908]=8'h00; mem['h5909]=8'h00; mem['h590A]=8'h00; mem['h590B]=8'h00;
    mem['h590C]=8'h00; mem['h590D]=8'h00; mem['h590E]=8'h00; mem['h590F]=8'h00;
    mem['h5910]=8'h00; mem['h5911]=8'h00; mem['h5912]=8'h00; mem['h5913]=8'h00;
    mem['h5914]=8'h00; mem['h5915]=8'h00; mem['h5916]=8'h00; mem['h5917]=8'h00;
    mem['h5918]=8'h00; mem['h5919]=8'h00; mem['h591A]=8'h00; mem['h591B]=8'h00;
    mem['h591C]=8'h00; mem['h591D]=8'h00; mem['h591E]=8'h00; mem['h591F]=8'h00;
    mem['h5920]=8'h00; mem['h5921]=8'h00; mem['h5922]=8'h00; mem['h5923]=8'h00;
    mem['h5924]=8'h00; mem['h5925]=8'h00; mem['h5926]=8'h00; mem['h5927]=8'h00;
    mem['h5928]=8'h00; mem['h5929]=8'h00; mem['h592A]=8'h00; mem['h592B]=8'h00;
    mem['h592C]=8'h00; mem['h592D]=8'h00; mem['h592E]=8'h00; mem['h592F]=8'h00;
    mem['h5930]=8'h00; mem['h5931]=8'h00; mem['h5932]=8'h00; mem['h5933]=8'h00;
    mem['h5934]=8'h00; mem['h5935]=8'h00; mem['h5936]=8'h00; mem['h5937]=8'h00;
    mem['h5938]=8'h00; mem['h5939]=8'h00; mem['h593A]=8'h00; mem['h593B]=8'h00;
    mem['h593C]=8'h00; mem['h593D]=8'h00; mem['h593E]=8'h00; mem['h593F]=8'h00;
    mem['h5940]=8'h00; mem['h5941]=8'h00; mem['h5942]=8'h00; mem['h5943]=8'h00;
    mem['h5944]=8'h00; mem['h5945]=8'h00; mem['h5946]=8'h00; mem['h5947]=8'h00;
    mem['h5948]=8'h00; mem['h5949]=8'h00; mem['h594A]=8'h00; mem['h594B]=8'h00;
    mem['h594C]=8'h00; mem['h594D]=8'h00; mem['h594E]=8'h00; mem['h594F]=8'h00;
    mem['h5950]=8'h00; mem['h5951]=8'h00; mem['h5952]=8'h00; mem['h5953]=8'h00;
    mem['h5954]=8'h00; mem['h5955]=8'h00; mem['h5956]=8'h00; mem['h5957]=8'h00;
    mem['h5958]=8'h00; mem['h5959]=8'h00; mem['h595A]=8'h00; mem['h595B]=8'h00;
    mem['h595C]=8'h00; mem['h595D]=8'h00; mem['h595E]=8'h00; mem['h595F]=8'h00;
    mem['h5960]=8'h00; mem['h5961]=8'h00; mem['h5962]=8'h00; mem['h5963]=8'h00;
    mem['h5964]=8'h00; mem['h5965]=8'h00; mem['h5966]=8'h00; mem['h5967]=8'h00;
    mem['h5968]=8'h00; mem['h5969]=8'h00; mem['h596A]=8'h00; mem['h596B]=8'h00;
    mem['h596C]=8'h00; mem['h596D]=8'h00; mem['h596E]=8'h00; mem['h596F]=8'h00;
    mem['h5970]=8'h00; mem['h5971]=8'h00; mem['h5972]=8'h00; mem['h5973]=8'h00;
    mem['h5974]=8'h00; mem['h5975]=8'h00; mem['h5976]=8'h00; mem['h5977]=8'h00;
    mem['h5978]=8'h00; mem['h5979]=8'h00; mem['h597A]=8'h00; mem['h597B]=8'h00;
    mem['h597C]=8'h00; mem['h597D]=8'h00; mem['h597E]=8'h00; mem['h597F]=8'h00;
    mem['h5980]=8'h00; mem['h5981]=8'h00; mem['h5982]=8'h00; mem['h5983]=8'h00;
    mem['h5984]=8'h00; mem['h5985]=8'h00; mem['h5986]=8'h00; mem['h5987]=8'h00;
    mem['h5988]=8'h00; mem['h5989]=8'h00; mem['h598A]=8'h00; mem['h598B]=8'h00;
    mem['h598C]=8'h00; mem['h598D]=8'h00; mem['h598E]=8'h00; mem['h598F]=8'h00;
    mem['h5990]=8'h00; mem['h5991]=8'h00; mem['h5992]=8'h00; mem['h5993]=8'h00;
    mem['h5994]=8'h00; mem['h5995]=8'h00; mem['h5996]=8'h00; mem['h5997]=8'h00;
    mem['h5998]=8'h00; mem['h5999]=8'h00; mem['h599A]=8'h00; mem['h599B]=8'h00;
    mem['h599C]=8'h00; mem['h599D]=8'h00; mem['h599E]=8'h00; mem['h599F]=8'h00;
    mem['h59A0]=8'h00; mem['h59A1]=8'h00; mem['h59A2]=8'h00; mem['h59A3]=8'h00;
    mem['h59A4]=8'h00; mem['h59A5]=8'h00; mem['h59A6]=8'h00; mem['h59A7]=8'h00;
    mem['h59A8]=8'h00; mem['h59A9]=8'h00; mem['h59AA]=8'h00; mem['h59AB]=8'h00;
    mem['h59AC]=8'h00; mem['h59AD]=8'h00; mem['h59AE]=8'h00; mem['h59AF]=8'h00;
    mem['h59B0]=8'h00; mem['h59B1]=8'h00; mem['h59B2]=8'h00; mem['h59B3]=8'h00;
    mem['h59B4]=8'h00; mem['h59B5]=8'h00; mem['h59B6]=8'h00; mem['h59B7]=8'h00;
    mem['h59B8]=8'h00; mem['h59B9]=8'h00; mem['h59BA]=8'h00; mem['h59BB]=8'h00;
    mem['h59BC]=8'h00; mem['h59BD]=8'h00; mem['h59BE]=8'h00; mem['h59BF]=8'h00;
    mem['h59C0]=8'h00; mem['h59C1]=8'h00; mem['h59C2]=8'h00; mem['h59C3]=8'h00;
    mem['h59C4]=8'h00; mem['h59C5]=8'h00; mem['h59C6]=8'h00; mem['h59C7]=8'h00;
    mem['h59C8]=8'h00; mem['h59C9]=8'h00; mem['h59CA]=8'h00; mem['h59CB]=8'h00;
    mem['h59CC]=8'h00; mem['h59CD]=8'h00; mem['h59CE]=8'h00; mem['h59CF]=8'h00;
    mem['h59D0]=8'h00; mem['h59D1]=8'h00; mem['h59D2]=8'h00; mem['h59D3]=8'h00;
    mem['h59D4]=8'h00; mem['h59D5]=8'h00; mem['h59D6]=8'h00; mem['h59D7]=8'h00;
    mem['h59D8]=8'h00; mem['h59D9]=8'h00; mem['h59DA]=8'h00; mem['h59DB]=8'h00;
    mem['h59DC]=8'h00; mem['h59DD]=8'h00; mem['h59DE]=8'h00; mem['h59DF]=8'h00;
    mem['h59E0]=8'h00; mem['h59E1]=8'h00; mem['h59E2]=8'h00; mem['h59E3]=8'h00;
    mem['h59E4]=8'h00; mem['h59E5]=8'h00; mem['h59E6]=8'h00; mem['h59E7]=8'h00;
    mem['h59E8]=8'h00; mem['h59E9]=8'h00; mem['h59EA]=8'h00; mem['h59EB]=8'h00;
    mem['h59EC]=8'h00; mem['h59ED]=8'h00; mem['h59EE]=8'h00; mem['h59EF]=8'h00;
    mem['h59F0]=8'h00; mem['h59F1]=8'h00; mem['h59F2]=8'h00; mem['h59F3]=8'h00;
    mem['h59F4]=8'h00; mem['h59F5]=8'h00; mem['h59F6]=8'h00; mem['h59F7]=8'h00;
    mem['h59F8]=8'h00; mem['h59F9]=8'h00; mem['h59FA]=8'h00; mem['h59FB]=8'h00;
    mem['h59FC]=8'h00; mem['h59FD]=8'h00; mem['h59FE]=8'h00; mem['h59FF]=8'h00;
    mem['h5A00]=8'h00; mem['h5A01]=8'h00; mem['h5A02]=8'h00; mem['h5A03]=8'h00;
    mem['h5A04]=8'h00; mem['h5A05]=8'h00; mem['h5A06]=8'h00; mem['h5A07]=8'h00;
    mem['h5A08]=8'h00; mem['h5A09]=8'h00; mem['h5A0A]=8'h00; mem['h5A0B]=8'h00;
    mem['h5A0C]=8'h00; mem['h5A0D]=8'h00; mem['h5A0E]=8'h00; mem['h5A0F]=8'h00;
    mem['h5A10]=8'h00; mem['h5A11]=8'h00; mem['h5A12]=8'h00; mem['h5A13]=8'h00;
    mem['h5A14]=8'h00; mem['h5A15]=8'h00; mem['h5A16]=8'h00; mem['h5A17]=8'h00;
    mem['h5A18]=8'h00; mem['h5A19]=8'h00; mem['h5A1A]=8'h00; mem['h5A1B]=8'h00;
    mem['h5A1C]=8'h00; mem['h5A1D]=8'h00; mem['h5A1E]=8'h00; mem['h5A1F]=8'h00;
    mem['h5A20]=8'h00; mem['h5A21]=8'h00; mem['h5A22]=8'h00; mem['h5A23]=8'h00;
    mem['h5A24]=8'h00; mem['h5A25]=8'h00; mem['h5A26]=8'h00; mem['h5A27]=8'h00;
    mem['h5A28]=8'h00; mem['h5A29]=8'h00; mem['h5A2A]=8'h00; mem['h5A2B]=8'h00;
    mem['h5A2C]=8'h00; mem['h5A2D]=8'h00; mem['h5A2E]=8'h00; mem['h5A2F]=8'h00;
    mem['h5A30]=8'h00; mem['h5A31]=8'h00; mem['h5A32]=8'h00; mem['h5A33]=8'h00;
    mem['h5A34]=8'h00; mem['h5A35]=8'h00; mem['h5A36]=8'h00; mem['h5A37]=8'h00;
    mem['h5A38]=8'h00; mem['h5A39]=8'h00; mem['h5A3A]=8'h00; mem['h5A3B]=8'h00;
    mem['h5A3C]=8'h00; mem['h5A3D]=8'h00; mem['h5A3E]=8'h00; mem['h5A3F]=8'h00;
    mem['h5A40]=8'h00; mem['h5A41]=8'h00; mem['h5A42]=8'h00; mem['h5A43]=8'h00;
    mem['h5A44]=8'h00; mem['h5A45]=8'h00; mem['h5A46]=8'h00; mem['h5A47]=8'h00;
    mem['h5A48]=8'h00; mem['h5A49]=8'h00; mem['h5A4A]=8'h00; mem['h5A4B]=8'h00;
    mem['h5A4C]=8'h00; mem['h5A4D]=8'h00; mem['h5A4E]=8'h00; mem['h5A4F]=8'h00;
    mem['h5A50]=8'h00; mem['h5A51]=8'h00; mem['h5A52]=8'h00; mem['h5A53]=8'h00;
    mem['h5A54]=8'h00; mem['h5A55]=8'h00; mem['h5A56]=8'h00; mem['h5A57]=8'h00;
    mem['h5A58]=8'h00; mem['h5A59]=8'h00; mem['h5A5A]=8'h00; mem['h5A5B]=8'h00;
    mem['h5A5C]=8'h00; mem['h5A5D]=8'h00; mem['h5A5E]=8'h00; mem['h5A5F]=8'h00;
    mem['h5A60]=8'h00; mem['h5A61]=8'h00; mem['h5A62]=8'h00; mem['h5A63]=8'h00;
    mem['h5A64]=8'h00; mem['h5A65]=8'h00; mem['h5A66]=8'h00; mem['h5A67]=8'h00;
    mem['h5A68]=8'h00; mem['h5A69]=8'h00; mem['h5A6A]=8'h00; mem['h5A6B]=8'h00;
    mem['h5A6C]=8'h00; mem['h5A6D]=8'h00; mem['h5A6E]=8'h00; mem['h5A6F]=8'h00;
    mem['h5A70]=8'h00; mem['h5A71]=8'h00; mem['h5A72]=8'h00; mem['h5A73]=8'h00;
    mem['h5A74]=8'h00; mem['h5A75]=8'h00; mem['h5A76]=8'h00; mem['h5A77]=8'h00;
    mem['h5A78]=8'h00; mem['h5A79]=8'h00; mem['h5A7A]=8'h00; mem['h5A7B]=8'h00;
    mem['h5A7C]=8'h00; mem['h5A7D]=8'h00; mem['h5A7E]=8'h00; mem['h5A7F]=8'h00;
    mem['h5A80]=8'h00; mem['h5A81]=8'h00; mem['h5A82]=8'h00; mem['h5A83]=8'h00;
    mem['h5A84]=8'h00; mem['h5A85]=8'h00; mem['h5A86]=8'h00; mem['h5A87]=8'h00;
    mem['h5A88]=8'h00; mem['h5A89]=8'h00; mem['h5A8A]=8'h00; mem['h5A8B]=8'h00;
    mem['h5A8C]=8'h00; mem['h5A8D]=8'h00; mem['h5A8E]=8'h00; mem['h5A8F]=8'h00;
    mem['h5A90]=8'h00; mem['h5A91]=8'h00; mem['h5A92]=8'h00; mem['h5A93]=8'h00;
    mem['h5A94]=8'h00; mem['h5A95]=8'h00; mem['h5A96]=8'h00; mem['h5A97]=8'h00;
    mem['h5A98]=8'h00; mem['h5A99]=8'h00; mem['h5A9A]=8'h00; mem['h5A9B]=8'h00;
    mem['h5A9C]=8'h00; mem['h5A9D]=8'h00; mem['h5A9E]=8'h00; mem['h5A9F]=8'h00;
    mem['h5AA0]=8'h00; mem['h5AA1]=8'h00; mem['h5AA2]=8'h00; mem['h5AA3]=8'h00;
    mem['h5AA4]=8'h00; mem['h5AA5]=8'h00; mem['h5AA6]=8'h00; mem['h5AA7]=8'h00;
    mem['h5AA8]=8'h00; mem['h5AA9]=8'h00; mem['h5AAA]=8'h00; mem['h5AAB]=8'h00;
    mem['h5AAC]=8'h00; mem['h5AAD]=8'h00; mem['h5AAE]=8'h00; mem['h5AAF]=8'h00;
    mem['h5AB0]=8'h00; mem['h5AB1]=8'h00; mem['h5AB2]=8'h00; mem['h5AB3]=8'h00;
    mem['h5AB4]=8'h00; mem['h5AB5]=8'h00; mem['h5AB6]=8'h00; mem['h5AB7]=8'h00;
    mem['h5AB8]=8'h00; mem['h5AB9]=8'h00; mem['h5ABA]=8'h00; mem['h5ABB]=8'h00;
    mem['h5ABC]=8'h00; mem['h5ABD]=8'h00; mem['h5ABE]=8'h00; mem['h5ABF]=8'h00;
    mem['h5AC0]=8'h00; mem['h5AC1]=8'h00; mem['h5AC2]=8'h00; mem['h5AC3]=8'h00;
    mem['h5AC4]=8'h00; mem['h5AC5]=8'h00; mem['h5AC6]=8'h00; mem['h5AC7]=8'h00;
    mem['h5AC8]=8'h00; mem['h5AC9]=8'h00; mem['h5ACA]=8'h00; mem['h5ACB]=8'h00;
    mem['h5ACC]=8'h00; mem['h5ACD]=8'h00; mem['h5ACE]=8'h00; mem['h5ACF]=8'h00;
    mem['h5AD0]=8'h00; mem['h5AD1]=8'h00; mem['h5AD2]=8'h00; mem['h5AD3]=8'h00;
    mem['h5AD4]=8'h00; mem['h5AD5]=8'h00; mem['h5AD6]=8'h00; mem['h5AD7]=8'h00;
    mem['h5AD8]=8'h00; mem['h5AD9]=8'h00; mem['h5ADA]=8'h00; mem['h5ADB]=8'h00;
    mem['h5ADC]=8'h00; mem['h5ADD]=8'h00; mem['h5ADE]=8'h00; mem['h5ADF]=8'h00;
    mem['h5AE0]=8'h00; mem['h5AE1]=8'h00; mem['h5AE2]=8'h00; mem['h5AE3]=8'h00;
    mem['h5AE4]=8'h00; mem['h5AE5]=8'h00; mem['h5AE6]=8'h00; mem['h5AE7]=8'h00;
    mem['h5AE8]=8'h00; mem['h5AE9]=8'h00; mem['h5AEA]=8'h00; mem['h5AEB]=8'h00;
    mem['h5AEC]=8'h00; mem['h5AED]=8'h00; mem['h5AEE]=8'h00; mem['h5AEF]=8'h00;
    mem['h5AF0]=8'h00; mem['h5AF1]=8'h00; mem['h5AF2]=8'h00; mem['h5AF3]=8'h00;
    mem['h5AF4]=8'h00; mem['h5AF5]=8'h00; mem['h5AF6]=8'h00; mem['h5AF7]=8'h00;
    mem['h5AF8]=8'h00; mem['h5AF9]=8'h00; mem['h5AFA]=8'h00; mem['h5AFB]=8'h00;
    mem['h5AFC]=8'h00; mem['h5AFD]=8'h00; mem['h5AFE]=8'h00; mem['h5AFF]=8'h00;
    mem['h5B00]=8'h00; mem['h5B01]=8'h00; mem['h5B02]=8'h00; mem['h5B03]=8'h00;
    mem['h5B04]=8'h00; mem['h5B05]=8'h00; mem['h5B06]=8'h00; mem['h5B07]=8'h00;
    mem['h5B08]=8'h00; mem['h5B09]=8'h00; mem['h5B0A]=8'h00; mem['h5B0B]=8'h00;
    mem['h5B0C]=8'h00; mem['h5B0D]=8'h00; mem['h5B0E]=8'h00; mem['h5B0F]=8'h00;
    mem['h5B10]=8'h00; mem['h5B11]=8'h00; mem['h5B12]=8'h00; mem['h5B13]=8'h00;
    mem['h5B14]=8'h00; mem['h5B15]=8'h00; mem['h5B16]=8'h00; mem['h5B17]=8'h00;
    mem['h5B18]=8'h00; mem['h5B19]=8'h00; mem['h5B1A]=8'h00; mem['h5B1B]=8'h00;
    mem['h5B1C]=8'h00; mem['h5B1D]=8'h00; mem['h5B1E]=8'h00; mem['h5B1F]=8'h00;
    mem['h5B20]=8'h00; mem['h5B21]=8'h00; mem['h5B22]=8'h00; mem['h5B23]=8'h00;
    mem['h5B24]=8'h00; mem['h5B25]=8'h00; mem['h5B26]=8'h00; mem['h5B27]=8'h00;
    mem['h5B28]=8'h00; mem['h5B29]=8'h00; mem['h5B2A]=8'h00; mem['h5B2B]=8'h00;
    mem['h5B2C]=8'h00; mem['h5B2D]=8'h00; mem['h5B2E]=8'h00; mem['h5B2F]=8'h00;
    mem['h5B30]=8'h00; mem['h5B31]=8'h00; mem['h5B32]=8'h00; mem['h5B33]=8'h00;
    mem['h5B34]=8'h00; mem['h5B35]=8'h00; mem['h5B36]=8'h00; mem['h5B37]=8'h00;
    mem['h5B38]=8'h00; mem['h5B39]=8'h00; mem['h5B3A]=8'h00; mem['h5B3B]=8'h00;
    mem['h5B3C]=8'h00; mem['h5B3D]=8'h00; mem['h5B3E]=8'h00; mem['h5B3F]=8'h00;
    mem['h5B40]=8'h00; mem['h5B41]=8'h00; mem['h5B42]=8'h00; mem['h5B43]=8'h00;
    mem['h5B44]=8'h00; mem['h5B45]=8'h00; mem['h5B46]=8'h00; mem['h5B47]=8'h00;
    mem['h5B48]=8'h00; mem['h5B49]=8'h00; mem['h5B4A]=8'h00; mem['h5B4B]=8'h00;
    mem['h5B4C]=8'h00; mem['h5B4D]=8'h00; mem['h5B4E]=8'h00; mem['h5B4F]=8'h00;
    mem['h5B50]=8'h00; mem['h5B51]=8'h00; mem['h5B52]=8'h00; mem['h5B53]=8'h00;
    mem['h5B54]=8'h00; mem['h5B55]=8'h00; mem['h5B56]=8'h00; mem['h5B57]=8'h00;
    mem['h5B58]=8'h00; mem['h5B59]=8'h00; mem['h5B5A]=8'h00; mem['h5B5B]=8'h00;
    mem['h5B5C]=8'h00; mem['h5B5D]=8'h00; mem['h5B5E]=8'h00; mem['h5B5F]=8'h00;
    mem['h5B60]=8'h00; mem['h5B61]=8'h00; mem['h5B62]=8'h00; mem['h5B63]=8'h00;
    mem['h5B64]=8'h00; mem['h5B65]=8'h00; mem['h5B66]=8'h00; mem['h5B67]=8'h00;
    mem['h5B68]=8'h00; mem['h5B69]=8'h00; mem['h5B6A]=8'h00; mem['h5B6B]=8'h00;
    mem['h5B6C]=8'h00; mem['h5B6D]=8'h00; mem['h5B6E]=8'h00; mem['h5B6F]=8'h00;
    mem['h5B70]=8'h00; mem['h5B71]=8'h00; mem['h5B72]=8'h00; mem['h5B73]=8'h00;
    mem['h5B74]=8'h00; mem['h5B75]=8'h00; mem['h5B76]=8'h00; mem['h5B77]=8'h00;
    mem['h5B78]=8'h00; mem['h5B79]=8'h00; mem['h5B7A]=8'h00; mem['h5B7B]=8'h00;
    mem['h5B7C]=8'h00; mem['h5B7D]=8'h00; mem['h5B7E]=8'h00; mem['h5B7F]=8'h00;
    mem['h5B80]=8'h00; mem['h5B81]=8'h00; mem['h5B82]=8'h00; mem['h5B83]=8'h00;
    mem['h5B84]=8'h00; mem['h5B85]=8'h00; mem['h5B86]=8'h00; mem['h5B87]=8'h00;
    mem['h5B88]=8'h00; mem['h5B89]=8'h00; mem['h5B8A]=8'h00; mem['h5B8B]=8'h00;
    mem['h5B8C]=8'h00; mem['h5B8D]=8'h00; mem['h5B8E]=8'h00; mem['h5B8F]=8'h00;
    mem['h5B90]=8'h00; mem['h5B91]=8'h00; mem['h5B92]=8'h00; mem['h5B93]=8'h00;
    mem['h5B94]=8'h00; mem['h5B95]=8'h00; mem['h5B96]=8'h00; mem['h5B97]=8'h00;
    mem['h5B98]=8'h00; mem['h5B99]=8'h00; mem['h5B9A]=8'h00; mem['h5B9B]=8'h00;
    mem['h5B9C]=8'h00; mem['h5B9D]=8'h00; mem['h5B9E]=8'h00; mem['h5B9F]=8'h00;
    mem['h5BA0]=8'h00; mem['h5BA1]=8'h00; mem['h5BA2]=8'h00; mem['h5BA3]=8'h00;
    mem['h5BA4]=8'h00; mem['h5BA5]=8'h00; mem['h5BA6]=8'h00; mem['h5BA7]=8'h00;
    mem['h5BA8]=8'h00; mem['h5BA9]=8'h00; mem['h5BAA]=8'h00; mem['h5BAB]=8'h00;
    mem['h5BAC]=8'h00; mem['h5BAD]=8'h00; mem['h5BAE]=8'h00; mem['h5BAF]=8'h00;
    mem['h5BB0]=8'h00; mem['h5BB1]=8'h00; mem['h5BB2]=8'h00; mem['h5BB3]=8'h00;
    mem['h5BB4]=8'h00; mem['h5BB5]=8'h00; mem['h5BB6]=8'h00; mem['h5BB7]=8'h00;
    mem['h5BB8]=8'h00; mem['h5BB9]=8'h00; mem['h5BBA]=8'h00; mem['h5BBB]=8'h00;
    mem['h5BBC]=8'h00; mem['h5BBD]=8'h00; mem['h5BBE]=8'h00; mem['h5BBF]=8'h00;
    mem['h5BC0]=8'h00; mem['h5BC1]=8'h00; mem['h5BC2]=8'h00; mem['h5BC3]=8'h00;
    mem['h5BC4]=8'h00; mem['h5BC5]=8'h00; mem['h5BC6]=8'h00; mem['h5BC7]=8'h00;
    mem['h5BC8]=8'h00; mem['h5BC9]=8'h00; mem['h5BCA]=8'h00; mem['h5BCB]=8'h00;
    mem['h5BCC]=8'h00; mem['h5BCD]=8'h00; mem['h5BCE]=8'h00; mem['h5BCF]=8'h00;
    mem['h5BD0]=8'h00; mem['h5BD1]=8'h00; mem['h5BD2]=8'h00; mem['h5BD3]=8'h00;
    mem['h5BD4]=8'h00; mem['h5BD5]=8'h00; mem['h5BD6]=8'h00; mem['h5BD7]=8'h00;
    mem['h5BD8]=8'h00; mem['h5BD9]=8'h00; mem['h5BDA]=8'h00; mem['h5BDB]=8'h00;
    mem['h5BDC]=8'h00; mem['h5BDD]=8'h00; mem['h5BDE]=8'h00; mem['h5BDF]=8'h00;
    mem['h5BE0]=8'h00; mem['h5BE1]=8'h00; mem['h5BE2]=8'h00; mem['h5BE3]=8'h00;
    mem['h5BE4]=8'h00; mem['h5BE5]=8'h00; mem['h5BE6]=8'h00; mem['h5BE7]=8'h00;
    mem['h5BE8]=8'h00; mem['h5BE9]=8'h00; mem['h5BEA]=8'h00; mem['h5BEB]=8'h00;
    mem['h5BEC]=8'h00; mem['h5BED]=8'h00; mem['h5BEE]=8'h00; mem['h5BEF]=8'h00;
    mem['h5BF0]=8'h00; mem['h5BF1]=8'h00; mem['h5BF2]=8'h00; mem['h5BF3]=8'h00;
    mem['h5BF4]=8'h00; mem['h5BF5]=8'h00; mem['h5BF6]=8'h00; mem['h5BF7]=8'h00;
    mem['h5BF8]=8'h00; mem['h5BF9]=8'h00; mem['h5BFA]=8'h00; mem['h5BFB]=8'h00;
    mem['h5BFC]=8'h00; mem['h5BFD]=8'h00; mem['h5BFE]=8'h00; mem['h5BFF]=8'h00;
    mem['h5C00]=8'h00; mem['h5C01]=8'h00; mem['h5C02]=8'h00; mem['h5C03]=8'h00;
    mem['h5C04]=8'h00; mem['h5C05]=8'h00; mem['h5C06]=8'h00; mem['h5C07]=8'h00;
    mem['h5C08]=8'h00; mem['h5C09]=8'h00; mem['h5C0A]=8'h00; mem['h5C0B]=8'h00;
    mem['h5C0C]=8'h00; mem['h5C0D]=8'h00; mem['h5C0E]=8'h00; mem['h5C0F]=8'h00;
    mem['h5C10]=8'h00; mem['h5C11]=8'h00; mem['h5C12]=8'h00; mem['h5C13]=8'h00;
    mem['h5C14]=8'h00; mem['h5C15]=8'h00; mem['h5C16]=8'h00; mem['h5C17]=8'h00;
    mem['h5C18]=8'h00; mem['h5C19]=8'h00; mem['h5C1A]=8'h00; mem['h5C1B]=8'h00;
    mem['h5C1C]=8'h00; mem['h5C1D]=8'h00; mem['h5C1E]=8'h00; mem['h5C1F]=8'h00;
    mem['h5C20]=8'h00; mem['h5C21]=8'h00; mem['h5C22]=8'h00; mem['h5C23]=8'h00;
    mem['h5C24]=8'h00; mem['h5C25]=8'h00; mem['h5C26]=8'h00; mem['h5C27]=8'h00;
    mem['h5C28]=8'h00; mem['h5C29]=8'h00; mem['h5C2A]=8'h00; mem['h5C2B]=8'h00;
    mem['h5C2C]=8'h00; mem['h5C2D]=8'h00; mem['h5C2E]=8'h00; mem['h5C2F]=8'h00;
    mem['h5C30]=8'h00; mem['h5C31]=8'h00; mem['h5C32]=8'h00; mem['h5C33]=8'h00;
    mem['h5C34]=8'h00; mem['h5C35]=8'h00; mem['h5C36]=8'h00; mem['h5C37]=8'h00;
    mem['h5C38]=8'h00; mem['h5C39]=8'h00; mem['h5C3A]=8'h00; mem['h5C3B]=8'h00;
    mem['h5C3C]=8'h00; mem['h5C3D]=8'h00; mem['h5C3E]=8'h00; mem['h5C3F]=8'h00;
    mem['h5C40]=8'h00; mem['h5C41]=8'h00; mem['h5C42]=8'h00; mem['h5C43]=8'h00;
    mem['h5C44]=8'h00; mem['h5C45]=8'h00; mem['h5C46]=8'h00; mem['h5C47]=8'h00;
    mem['h5C48]=8'h00; mem['h5C49]=8'h00; mem['h5C4A]=8'h00; mem['h5C4B]=8'h00;
    mem['h5C4C]=8'h00; mem['h5C4D]=8'h00; mem['h5C4E]=8'h00; mem['h5C4F]=8'h00;
    mem['h5C50]=8'h00; mem['h5C51]=8'h00; mem['h5C52]=8'h00; mem['h5C53]=8'h00;
    mem['h5C54]=8'h00; mem['h5C55]=8'h00; mem['h5C56]=8'h00; mem['h5C57]=8'h00;
    mem['h5C58]=8'h00; mem['h5C59]=8'h00; mem['h5C5A]=8'h00; mem['h5C5B]=8'h00;
    mem['h5C5C]=8'h00; mem['h5C5D]=8'h00; mem['h5C5E]=8'h00; mem['h5C5F]=8'h00;
    mem['h5C60]=8'h00; mem['h5C61]=8'h00; mem['h5C62]=8'h00; mem['h5C63]=8'h00;
    mem['h5C64]=8'h00; mem['h5C65]=8'h00; mem['h5C66]=8'h00; mem['h5C67]=8'h00;
    mem['h5C68]=8'h00; mem['h5C69]=8'h00; mem['h5C6A]=8'h00; mem['h5C6B]=8'h00;
    mem['h5C6C]=8'h00; mem['h5C6D]=8'h00; mem['h5C6E]=8'h00; mem['h5C6F]=8'h00;
    mem['h5C70]=8'h00; mem['h5C71]=8'h00; mem['h5C72]=8'h00; mem['h5C73]=8'h00;
    mem['h5C74]=8'h00; mem['h5C75]=8'h00; mem['h5C76]=8'h00; mem['h5C77]=8'h00;
    mem['h5C78]=8'h00; mem['h5C79]=8'h00; mem['h5C7A]=8'h00; mem['h5C7B]=8'h00;
    mem['h5C7C]=8'h00; mem['h5C7D]=8'h00; mem['h5C7E]=8'h00; mem['h5C7F]=8'h00;
    mem['h5C80]=8'h00; mem['h5C81]=8'h00; mem['h5C82]=8'h00; mem['h5C83]=8'h00;
    mem['h5C84]=8'h00; mem['h5C85]=8'h00; mem['h5C86]=8'h00; mem['h5C87]=8'h00;
    mem['h5C88]=8'h00; mem['h5C89]=8'h00; mem['h5C8A]=8'h00; mem['h5C8B]=8'h00;
    mem['h5C8C]=8'h00; mem['h5C8D]=8'h00; mem['h5C8E]=8'h00; mem['h5C8F]=8'h00;
    mem['h5C90]=8'h00; mem['h5C91]=8'h00; mem['h5C92]=8'h00; mem['h5C93]=8'h00;
    mem['h5C94]=8'h00; mem['h5C95]=8'h00; mem['h5C96]=8'h00; mem['h5C97]=8'h00;
    mem['h5C98]=8'h00; mem['h5C99]=8'h00; mem['h5C9A]=8'h00; mem['h5C9B]=8'h00;
    mem['h5C9C]=8'h00; mem['h5C9D]=8'h00; mem['h5C9E]=8'h00; mem['h5C9F]=8'h00;
    mem['h5CA0]=8'h00; mem['h5CA1]=8'h00; mem['h5CA2]=8'h00; mem['h5CA3]=8'h00;
    mem['h5CA4]=8'h00; mem['h5CA5]=8'h00; mem['h5CA6]=8'h00; mem['h5CA7]=8'h00;
    mem['h5CA8]=8'h00; mem['h5CA9]=8'h00; mem['h5CAA]=8'h00; mem['h5CAB]=8'h00;
    mem['h5CAC]=8'h00; mem['h5CAD]=8'h00; mem['h5CAE]=8'h00; mem['h5CAF]=8'h00;
    mem['h5CB0]=8'h00; mem['h5CB1]=8'h00; mem['h5CB2]=8'h00; mem['h5CB3]=8'h00;
    mem['h5CB4]=8'h00; mem['h5CB5]=8'h00; mem['h5CB6]=8'h00; mem['h5CB7]=8'h00;
    mem['h5CB8]=8'h00; mem['h5CB9]=8'h00; mem['h5CBA]=8'h00; mem['h5CBB]=8'h00;
    mem['h5CBC]=8'h00; mem['h5CBD]=8'h00; mem['h5CBE]=8'h00; mem['h5CBF]=8'h00;
    mem['h5CC0]=8'h00; mem['h5CC1]=8'h00; mem['h5CC2]=8'h00; mem['h5CC3]=8'h00;
    mem['h5CC4]=8'h00; mem['h5CC5]=8'h00; mem['h5CC6]=8'h00; mem['h5CC7]=8'h00;
    mem['h5CC8]=8'h00; mem['h5CC9]=8'h00; mem['h5CCA]=8'h00; mem['h5CCB]=8'h00;
    mem['h5CCC]=8'h00; mem['h5CCD]=8'h00; mem['h5CCE]=8'h00; mem['h5CCF]=8'h00;
    mem['h5CD0]=8'h00; mem['h5CD1]=8'h00; mem['h5CD2]=8'h00; mem['h5CD3]=8'h00;
    mem['h5CD4]=8'h00; mem['h5CD5]=8'h00; mem['h5CD6]=8'h00; mem['h5CD7]=8'h00;
    mem['h5CD8]=8'h00; mem['h5CD9]=8'h00; mem['h5CDA]=8'h00; mem['h5CDB]=8'h00;
    mem['h5CDC]=8'h00; mem['h5CDD]=8'h00; mem['h5CDE]=8'h00; mem['h5CDF]=8'h00;
    mem['h5CE0]=8'h00; mem['h5CE1]=8'h00; mem['h5CE2]=8'h00; mem['h5CE3]=8'h00;
    mem['h5CE4]=8'h00; mem['h5CE5]=8'h00; mem['h5CE6]=8'h00; mem['h5CE7]=8'h00;
    mem['h5CE8]=8'h00; mem['h5CE9]=8'h00; mem['h5CEA]=8'h00; mem['h5CEB]=8'h00;
    mem['h5CEC]=8'h00; mem['h5CED]=8'h00; mem['h5CEE]=8'h00; mem['h5CEF]=8'h00;
    mem['h5CF0]=8'h00; mem['h5CF1]=8'h00; mem['h5CF2]=8'h00; mem['h5CF3]=8'h00;
    mem['h5CF4]=8'h00; mem['h5CF5]=8'h00; mem['h5CF6]=8'h00; mem['h5CF7]=8'h00;
    mem['h5CF8]=8'h00; mem['h5CF9]=8'h00; mem['h5CFA]=8'h00; mem['h5CFB]=8'h00;
    mem['h5CFC]=8'h00; mem['h5CFD]=8'h00; mem['h5CFE]=8'h00; mem['h5CFF]=8'h00;
    mem['h5D00]=8'h00; mem['h5D01]=8'h00; mem['h5D02]=8'h00; mem['h5D03]=8'h00;
    mem['h5D04]=8'h00; mem['h5D05]=8'h00; mem['h5D06]=8'h00; mem['h5D07]=8'h00;
    mem['h5D08]=8'h00; mem['h5D09]=8'h00; mem['h5D0A]=8'h00; mem['h5D0B]=8'h00;
    mem['h5D0C]=8'h00; mem['h5D0D]=8'h00; mem['h5D0E]=8'h00; mem['h5D0F]=8'h00;
    mem['h5D10]=8'h00; mem['h5D11]=8'h00; mem['h5D12]=8'h00; mem['h5D13]=8'h00;
    mem['h5D14]=8'h00; mem['h5D15]=8'h00; mem['h5D16]=8'h00; mem['h5D17]=8'h00;
    mem['h5D18]=8'h00; mem['h5D19]=8'h00; mem['h5D1A]=8'h00; mem['h5D1B]=8'h00;
    mem['h5D1C]=8'h00; mem['h5D1D]=8'h00; mem['h5D1E]=8'h00; mem['h5D1F]=8'h00;
    mem['h5D20]=8'h00; mem['h5D21]=8'h00; mem['h5D22]=8'h00; mem['h5D23]=8'h00;
    mem['h5D24]=8'h00; mem['h5D25]=8'h00; mem['h5D26]=8'h00; mem['h5D27]=8'h00;
    mem['h5D28]=8'h00; mem['h5D29]=8'h00; mem['h5D2A]=8'h00; mem['h5D2B]=8'h00;
    mem['h5D2C]=8'h00; mem['h5D2D]=8'h00; mem['h5D2E]=8'h00; mem['h5D2F]=8'h00;
    mem['h5D30]=8'h00; mem['h5D31]=8'h00; mem['h5D32]=8'h00; mem['h5D33]=8'h00;
    mem['h5D34]=8'h00; mem['h5D35]=8'h00; mem['h5D36]=8'h00; mem['h5D37]=8'h00;
    mem['h5D38]=8'h00; mem['h5D39]=8'h00; mem['h5D3A]=8'h00; mem['h5D3B]=8'h00;
    mem['h5D3C]=8'h00; mem['h5D3D]=8'h00; mem['h5D3E]=8'h00; mem['h5D3F]=8'h00;
    mem['h5D40]=8'h00; mem['h5D41]=8'h00; mem['h5D42]=8'h00; mem['h5D43]=8'h00;
    mem['h5D44]=8'h00; mem['h5D45]=8'h00; mem['h5D46]=8'h00; mem['h5D47]=8'h00;
    mem['h5D48]=8'h00; mem['h5D49]=8'h00; mem['h5D4A]=8'h00; mem['h5D4B]=8'h00;
    mem['h5D4C]=8'h00; mem['h5D4D]=8'h00; mem['h5D4E]=8'h00; mem['h5D4F]=8'h00;
    mem['h5D50]=8'h00; mem['h5D51]=8'h00; mem['h5D52]=8'h00; mem['h5D53]=8'h00;
    mem['h5D54]=8'h00; mem['h5D55]=8'h00; mem['h5D56]=8'h00; mem['h5D57]=8'h00;
    mem['h5D58]=8'h00; mem['h5D59]=8'h00; mem['h5D5A]=8'h00; mem['h5D5B]=8'h00;
    mem['h5D5C]=8'h00; mem['h5D5D]=8'h00; mem['h5D5E]=8'h00; mem['h5D5F]=8'h00;
    mem['h5D60]=8'h00; mem['h5D61]=8'h00; mem['h5D62]=8'h00; mem['h5D63]=8'h00;
    mem['h5D64]=8'h00; mem['h5D65]=8'h00; mem['h5D66]=8'h00; mem['h5D67]=8'h00;
    mem['h5D68]=8'h00; mem['h5D69]=8'h00; mem['h5D6A]=8'h00; mem['h5D6B]=8'h00;
    mem['h5D6C]=8'h00; mem['h5D6D]=8'h00; mem['h5D6E]=8'h00; mem['h5D6F]=8'h00;
    mem['h5D70]=8'h00; mem['h5D71]=8'h00; mem['h5D72]=8'h00; mem['h5D73]=8'h00;
    mem['h5D74]=8'h00; mem['h5D75]=8'h00; mem['h5D76]=8'h00; mem['h5D77]=8'h00;
    mem['h5D78]=8'h00; mem['h5D79]=8'h00; mem['h5D7A]=8'h00; mem['h5D7B]=8'h00;
    mem['h5D7C]=8'h00; mem['h5D7D]=8'h00; mem['h5D7E]=8'h00; mem['h5D7F]=8'h00;
    mem['h5D80]=8'h00; mem['h5D81]=8'h00; mem['h5D82]=8'h00; mem['h5D83]=8'h00;
    mem['h5D84]=8'h00; mem['h5D85]=8'h00; mem['h5D86]=8'h00; mem['h5D87]=8'h00;
    mem['h5D88]=8'h00; mem['h5D89]=8'h00; mem['h5D8A]=8'h00; mem['h5D8B]=8'h00;
    mem['h5D8C]=8'h00; mem['h5D8D]=8'h00; mem['h5D8E]=8'h00; mem['h5D8F]=8'h00;
    mem['h5D90]=8'h00; mem['h5D91]=8'h00; mem['h5D92]=8'h00; mem['h5D93]=8'h00;
    mem['h5D94]=8'h00; mem['h5D95]=8'h00; mem['h5D96]=8'h00; mem['h5D97]=8'h00;
    mem['h5D98]=8'h00; mem['h5D99]=8'h00; mem['h5D9A]=8'h00; mem['h5D9B]=8'h00;
    mem['h5D9C]=8'h00; mem['h5D9D]=8'h00; mem['h5D9E]=8'h00; mem['h5D9F]=8'h00;
    mem['h5DA0]=8'h00; mem['h5DA1]=8'h00; mem['h5DA2]=8'h00; mem['h5DA3]=8'h00;
    mem['h5DA4]=8'h00; mem['h5DA5]=8'h00; mem['h5DA6]=8'h00; mem['h5DA7]=8'h00;
    mem['h5DA8]=8'h00; mem['h5DA9]=8'h00; mem['h5DAA]=8'h00; mem['h5DAB]=8'h00;
    mem['h5DAC]=8'h00; mem['h5DAD]=8'h00; mem['h5DAE]=8'h00; mem['h5DAF]=8'h00;
    mem['h5DB0]=8'h00; mem['h5DB1]=8'h00; mem['h5DB2]=8'h00; mem['h5DB3]=8'h00;
    mem['h5DB4]=8'h00; mem['h5DB5]=8'h00; mem['h5DB6]=8'h00; mem['h5DB7]=8'h00;
    mem['h5DB8]=8'h00; mem['h5DB9]=8'h00; mem['h5DBA]=8'h00; mem['h5DBB]=8'h00;
    mem['h5DBC]=8'h00; mem['h5DBD]=8'h00; mem['h5DBE]=8'h00; mem['h5DBF]=8'h00;
    mem['h5DC0]=8'h00; mem['h5DC1]=8'h00; mem['h5DC2]=8'h00; mem['h5DC3]=8'h00;
    mem['h5DC4]=8'h00; mem['h5DC5]=8'h00; mem['h5DC6]=8'h00; mem['h5DC7]=8'h00;
    mem['h5DC8]=8'h00; mem['h5DC9]=8'h00; mem['h5DCA]=8'h00; mem['h5DCB]=8'h00;
    mem['h5DCC]=8'h00; mem['h5DCD]=8'h00; mem['h5DCE]=8'h00; mem['h5DCF]=8'h00;
    mem['h5DD0]=8'h00; mem['h5DD1]=8'h00; mem['h5DD2]=8'h00; mem['h5DD3]=8'h00;
    mem['h5DD4]=8'h00; mem['h5DD5]=8'h00; mem['h5DD6]=8'h00; mem['h5DD7]=8'h00;
    mem['h5DD8]=8'h00; mem['h5DD9]=8'h00; mem['h5DDA]=8'h00; mem['h5DDB]=8'h00;
    mem['h5DDC]=8'h00; mem['h5DDD]=8'h00; mem['h5DDE]=8'h00; mem['h5DDF]=8'h00;
    mem['h5DE0]=8'h00; mem['h5DE1]=8'h00; mem['h5DE2]=8'h00; mem['h5DE3]=8'h00;
    mem['h5DE4]=8'h00; mem['h5DE5]=8'h00; mem['h5DE6]=8'h00; mem['h5DE7]=8'h00;
    mem['h5DE8]=8'h00; mem['h5DE9]=8'h00; mem['h5DEA]=8'h00; mem['h5DEB]=8'h00;
    mem['h5DEC]=8'h00; mem['h5DED]=8'h00; mem['h5DEE]=8'h00; mem['h5DEF]=8'h00;
    mem['h5DF0]=8'h00; mem['h5DF1]=8'h00; mem['h5DF2]=8'h00; mem['h5DF3]=8'h00;
    mem['h5DF4]=8'h00; mem['h5DF5]=8'h00; mem['h5DF6]=8'h00; mem['h5DF7]=8'h00;
    mem['h5DF8]=8'h00; mem['h5DF9]=8'h00; mem['h5DFA]=8'h00; mem['h5DFB]=8'h00;
    mem['h5DFC]=8'h00; mem['h5DFD]=8'h00; mem['h5DFE]=8'h00; mem['h5DFF]=8'h00;
    mem['h5E00]=8'h00; mem['h5E01]=8'h00; mem['h5E02]=8'h00; mem['h5E03]=8'h00;
    mem['h5E04]=8'h00; mem['h5E05]=8'h00; mem['h5E06]=8'h00; mem['h5E07]=8'h00;
    mem['h5E08]=8'h00; mem['h5E09]=8'h00; mem['h5E0A]=8'h00; mem['h5E0B]=8'h00;
    mem['h5E0C]=8'h00; mem['h5E0D]=8'h00; mem['h5E0E]=8'h00; mem['h5E0F]=8'h00;
    mem['h5E10]=8'h00; mem['h5E11]=8'h00; mem['h5E12]=8'h00; mem['h5E13]=8'h00;
    mem['h5E14]=8'h00; mem['h5E15]=8'h00; mem['h5E16]=8'h00; mem['h5E17]=8'h00;
    mem['h5E18]=8'h00; mem['h5E19]=8'h00; mem['h5E1A]=8'h00; mem['h5E1B]=8'h00;
    mem['h5E1C]=8'h00; mem['h5E1D]=8'h00; mem['h5E1E]=8'h00; mem['h5E1F]=8'h00;
    mem['h5E20]=8'h00; mem['h5E21]=8'h00; mem['h5E22]=8'h00; mem['h5E23]=8'h00;
    mem['h5E24]=8'h00; mem['h5E25]=8'h00; mem['h5E26]=8'h00; mem['h5E27]=8'h00;
    mem['h5E28]=8'h00; mem['h5E29]=8'h00; mem['h5E2A]=8'h00; mem['h5E2B]=8'h00;
    mem['h5E2C]=8'h00; mem['h5E2D]=8'h00; mem['h5E2E]=8'h00; mem['h5E2F]=8'h00;
    mem['h5E30]=8'h00; mem['h5E31]=8'h00; mem['h5E32]=8'h00; mem['h5E33]=8'h00;
    mem['h5E34]=8'h00; mem['h5E35]=8'h00; mem['h5E36]=8'h00; mem['h5E37]=8'h00;
    mem['h5E38]=8'h00; mem['h5E39]=8'h00; mem['h5E3A]=8'h00; mem['h5E3B]=8'h00;
    mem['h5E3C]=8'h00; mem['h5E3D]=8'h00; mem['h5E3E]=8'h00; mem['h5E3F]=8'h00;
    mem['h5E40]=8'h00; mem['h5E41]=8'h00; mem['h5E42]=8'h00; mem['h5E43]=8'h00;
    mem['h5E44]=8'h00; mem['h5E45]=8'h00; mem['h5E46]=8'h00; mem['h5E47]=8'h00;
    mem['h5E48]=8'h00; mem['h5E49]=8'h00; mem['h5E4A]=8'h00; mem['h5E4B]=8'h00;
    mem['h5E4C]=8'h00; mem['h5E4D]=8'h00; mem['h5E4E]=8'h00; mem['h5E4F]=8'h00;
    mem['h5E50]=8'h00; mem['h5E51]=8'h00; mem['h5E52]=8'h00; mem['h5E53]=8'h00;
    mem['h5E54]=8'h00; mem['h5E55]=8'h00; mem['h5E56]=8'h00; mem['h5E57]=8'h00;
    mem['h5E58]=8'h00; mem['h5E59]=8'h00; mem['h5E5A]=8'h00; mem['h5E5B]=8'h00;
    mem['h5E5C]=8'h00; mem['h5E5D]=8'h00; mem['h5E5E]=8'h00; mem['h5E5F]=8'h00;
    mem['h5E60]=8'h00; mem['h5E61]=8'h00; mem['h5E62]=8'h00; mem['h5E63]=8'h00;
    mem['h5E64]=8'h00; mem['h5E65]=8'h00; mem['h5E66]=8'h00; mem['h5E67]=8'h00;
    mem['h5E68]=8'h00; mem['h5E69]=8'h00; mem['h5E6A]=8'h00; mem['h5E6B]=8'h00;
    mem['h5E6C]=8'h00; mem['h5E6D]=8'h00; mem['h5E6E]=8'h00; mem['h5E6F]=8'h00;
    mem['h5E70]=8'h00; mem['h5E71]=8'h00; mem['h5E72]=8'h00; mem['h5E73]=8'h00;
    mem['h5E74]=8'h00; mem['h5E75]=8'h00; mem['h5E76]=8'h00; mem['h5E77]=8'h00;
    mem['h5E78]=8'h00; mem['h5E79]=8'h00; mem['h5E7A]=8'h00; mem['h5E7B]=8'h00;
    mem['h5E7C]=8'h00; mem['h5E7D]=8'h00; mem['h5E7E]=8'h00; mem['h5E7F]=8'h00;
    mem['h5E80]=8'h00; mem['h5E81]=8'h00; mem['h5E82]=8'h00; mem['h5E83]=8'h00;
    mem['h5E84]=8'h00; mem['h5E85]=8'h00; mem['h5E86]=8'h00; mem['h5E87]=8'h00;
    mem['h5E88]=8'h00; mem['h5E89]=8'h00; mem['h5E8A]=8'h00; mem['h5E8B]=8'h00;
    mem['h5E8C]=8'h00; mem['h5E8D]=8'h00; mem['h5E8E]=8'h00; mem['h5E8F]=8'h00;
    mem['h5E90]=8'h00; mem['h5E91]=8'h00; mem['h5E92]=8'h00; mem['h5E93]=8'h00;
    mem['h5E94]=8'h00; mem['h5E95]=8'h00; mem['h5E96]=8'h00; mem['h5E97]=8'h00;
    mem['h5E98]=8'h00; mem['h5E99]=8'h00; mem['h5E9A]=8'h00; mem['h5E9B]=8'h00;
    mem['h5E9C]=8'h00; mem['h5E9D]=8'h00; mem['h5E9E]=8'h00; mem['h5E9F]=8'h00;
    mem['h5EA0]=8'h00; mem['h5EA1]=8'h00; mem['h5EA2]=8'h00; mem['h5EA3]=8'h00;
    mem['h5EA4]=8'h00; mem['h5EA5]=8'h00; mem['h5EA6]=8'h00; mem['h5EA7]=8'h00;
    mem['h5EA8]=8'h00; mem['h5EA9]=8'h00; mem['h5EAA]=8'h00; mem['h5EAB]=8'h00;
    mem['h5EAC]=8'h00; mem['h5EAD]=8'h00; mem['h5EAE]=8'h00; mem['h5EAF]=8'h00;
    mem['h5EB0]=8'h00; mem['h5EB1]=8'h00; mem['h5EB2]=8'h00; mem['h5EB3]=8'h00;
    mem['h5EB4]=8'h00; mem['h5EB5]=8'h00; mem['h5EB6]=8'h00; mem['h5EB7]=8'h00;
    mem['h5EB8]=8'h00; mem['h5EB9]=8'h00; mem['h5EBA]=8'h00; mem['h5EBB]=8'h00;
    mem['h5EBC]=8'h00; mem['h5EBD]=8'h00; mem['h5EBE]=8'h00; mem['h5EBF]=8'h00;
    mem['h5EC0]=8'h00; mem['h5EC1]=8'h00; mem['h5EC2]=8'h00; mem['h5EC3]=8'h00;
    mem['h5EC4]=8'h00; mem['h5EC5]=8'h00; mem['h5EC6]=8'h00; mem['h5EC7]=8'h00;
    mem['h5EC8]=8'h00; mem['h5EC9]=8'h00; mem['h5ECA]=8'h00; mem['h5ECB]=8'h00;
    mem['h5ECC]=8'h00; mem['h5ECD]=8'h00; mem['h5ECE]=8'h00; mem['h5ECF]=8'h00;
    mem['h5ED0]=8'h00; mem['h5ED1]=8'h00; mem['h5ED2]=8'h00; mem['h5ED3]=8'h00;
    mem['h5ED4]=8'h00; mem['h5ED5]=8'h00; mem['h5ED6]=8'h00; mem['h5ED7]=8'h00;
    mem['h5ED8]=8'h00; mem['h5ED9]=8'h00; mem['h5EDA]=8'h00; mem['h5EDB]=8'h00;
    mem['h5EDC]=8'h00; mem['h5EDD]=8'h00; mem['h5EDE]=8'h00; mem['h5EDF]=8'h00;
    mem['h5EE0]=8'h00; mem['h5EE1]=8'h00; mem['h5EE2]=8'h00; mem['h5EE3]=8'h00;
    mem['h5EE4]=8'h00; mem['h5EE5]=8'h00; mem['h5EE6]=8'h00; mem['h5EE7]=8'h00;
    mem['h5EE8]=8'h00; mem['h5EE9]=8'h00; mem['h5EEA]=8'h00; mem['h5EEB]=8'h00;
    mem['h5EEC]=8'h00; mem['h5EED]=8'h00; mem['h5EEE]=8'h00; mem['h5EEF]=8'h00;
    mem['h5EF0]=8'h00; mem['h5EF1]=8'h00; mem['h5EF2]=8'h00; mem['h5EF3]=8'h00;
    mem['h5EF4]=8'h00; mem['h5EF5]=8'h00; mem['h5EF6]=8'h00; mem['h5EF7]=8'h00;
    mem['h5EF8]=8'h00; mem['h5EF9]=8'h00; mem['h5EFA]=8'h00; mem['h5EFB]=8'h00;
    mem['h5EFC]=8'h00; mem['h5EFD]=8'h00; mem['h5EFE]=8'h00; mem['h5EFF]=8'h00;
    mem['h5F00]=8'h00; mem['h5F01]=8'h00; mem['h5F02]=8'h00; mem['h5F03]=8'h00;
    mem['h5F04]=8'h00; mem['h5F05]=8'h00; mem['h5F06]=8'h00; mem['h5F07]=8'h00;
    mem['h5F08]=8'h00; mem['h5F09]=8'h00; mem['h5F0A]=8'h00; mem['h5F0B]=8'h00;
    mem['h5F0C]=8'h00; mem['h5F0D]=8'h00; mem['h5F0E]=8'h00; mem['h5F0F]=8'h00;
    mem['h5F10]=8'h00; mem['h5F11]=8'h00; mem['h5F12]=8'h00; mem['h5F13]=8'h00;
    mem['h5F14]=8'h00; mem['h5F15]=8'h00; mem['h5F16]=8'h00; mem['h5F17]=8'h00;
    mem['h5F18]=8'h00; mem['h5F19]=8'h00; mem['h5F1A]=8'h00; mem['h5F1B]=8'h00;
    mem['h5F1C]=8'h00; mem['h5F1D]=8'h00; mem['h5F1E]=8'h00; mem['h5F1F]=8'h00;
    mem['h5F20]=8'h00; mem['h5F21]=8'h00; mem['h5F22]=8'h00; mem['h5F23]=8'h00;
    mem['h5F24]=8'h00; mem['h5F25]=8'h00; mem['h5F26]=8'h00; mem['h5F27]=8'h00;
    mem['h5F28]=8'h00; mem['h5F29]=8'h00; mem['h5F2A]=8'h00; mem['h5F2B]=8'h00;
    mem['h5F2C]=8'h00; mem['h5F2D]=8'h00; mem['h5F2E]=8'h00; mem['h5F2F]=8'h00;
    mem['h5F30]=8'h00; mem['h5F31]=8'h00; mem['h5F32]=8'h00; mem['h5F33]=8'h00;
    mem['h5F34]=8'h00; mem['h5F35]=8'h00; mem['h5F36]=8'h00; mem['h5F37]=8'h00;
    mem['h5F38]=8'h00; mem['h5F39]=8'h00; mem['h5F3A]=8'h00; mem['h5F3B]=8'h00;
    mem['h5F3C]=8'h00; mem['h5F3D]=8'h00; mem['h5F3E]=8'h00; mem['h5F3F]=8'h00;
    mem['h5F40]=8'h00; mem['h5F41]=8'h00; mem['h5F42]=8'h00; mem['h5F43]=8'h00;
    mem['h5F44]=8'h00; mem['h5F45]=8'h00; mem['h5F46]=8'h00; mem['h5F47]=8'h00;
    mem['h5F48]=8'h00; mem['h5F49]=8'h00; mem['h5F4A]=8'h00; mem['h5F4B]=8'h00;
    mem['h5F4C]=8'h00; mem['h5F4D]=8'h00; mem['h5F4E]=8'h00; mem['h5F4F]=8'h00;
    mem['h5F50]=8'h00; mem['h5F51]=8'h00; mem['h5F52]=8'h00; mem['h5F53]=8'h00;
    mem['h5F54]=8'h00; mem['h5F55]=8'h00; mem['h5F56]=8'h00; mem['h5F57]=8'h00;
    mem['h5F58]=8'h00; mem['h5F59]=8'h00; mem['h5F5A]=8'h00; mem['h5F5B]=8'h00;
    mem['h5F5C]=8'h00; mem['h5F5D]=8'h00; mem['h5F5E]=8'h00; mem['h5F5F]=8'h00;
    mem['h5F60]=8'h00; mem['h5F61]=8'h00; mem['h5F62]=8'h00; mem['h5F63]=8'h00;
    mem['h5F64]=8'h00; mem['h5F65]=8'h00; mem['h5F66]=8'h00; mem['h5F67]=8'h00;
    mem['h5F68]=8'h00; mem['h5F69]=8'h00; mem['h5F6A]=8'h00; mem['h5F6B]=8'h00;
    mem['h5F6C]=8'h00; mem['h5F6D]=8'h00; mem['h5F6E]=8'h00; mem['h5F6F]=8'h00;
    mem['h5F70]=8'h00; mem['h5F71]=8'h00; mem['h5F72]=8'h00; mem['h5F73]=8'h00;
    mem['h5F74]=8'h00; mem['h5F75]=8'h00; mem['h5F76]=8'h00; mem['h5F77]=8'h00;
    mem['h5F78]=8'h00; mem['h5F79]=8'h00; mem['h5F7A]=8'h00; mem['h5F7B]=8'h00;
    mem['h5F7C]=8'h00; mem['h5F7D]=8'h00; mem['h5F7E]=8'h00; mem['h5F7F]=8'h00;
    mem['h5F80]=8'h00; mem['h5F81]=8'h00; mem['h5F82]=8'h00; mem['h5F83]=8'h00;
    mem['h5F84]=8'h00; mem['h5F85]=8'h00; mem['h5F86]=8'h00; mem['h5F87]=8'h00;
    mem['h5F88]=8'h00; mem['h5F89]=8'h00; mem['h5F8A]=8'h00; mem['h5F8B]=8'h00;
    mem['h5F8C]=8'h00; mem['h5F8D]=8'h00; mem['h5F8E]=8'h00; mem['h5F8F]=8'h00;
    mem['h5F90]=8'h00; mem['h5F91]=8'h00; mem['h5F92]=8'h00; mem['h5F93]=8'h00;
    mem['h5F94]=8'h00; mem['h5F95]=8'h00; mem['h5F96]=8'h00; mem['h5F97]=8'h00;
    mem['h5F98]=8'h00; mem['h5F99]=8'h00; mem['h5F9A]=8'h00; mem['h5F9B]=8'h00;
    mem['h5F9C]=8'h00; mem['h5F9D]=8'h00; mem['h5F9E]=8'h00; mem['h5F9F]=8'h00;
    mem['h5FA0]=8'h00; mem['h5FA1]=8'h00; mem['h5FA2]=8'h00; mem['h5FA3]=8'h00;
    mem['h5FA4]=8'h00; mem['h5FA5]=8'h00; mem['h5FA6]=8'h00; mem['h5FA7]=8'h00;
    mem['h5FA8]=8'h00; mem['h5FA9]=8'h00; mem['h5FAA]=8'h00; mem['h5FAB]=8'h00;
    mem['h5FAC]=8'h00; mem['h5FAD]=8'h00; mem['h5FAE]=8'h00; mem['h5FAF]=8'h00;
    mem['h5FB0]=8'h00; mem['h5FB1]=8'h00; mem['h5FB2]=8'h00; mem['h5FB3]=8'h00;
    mem['h5FB4]=8'h00; mem['h5FB5]=8'h00; mem['h5FB6]=8'h00; mem['h5FB7]=8'h00;
    mem['h5FB8]=8'h00; mem['h5FB9]=8'h00; mem['h5FBA]=8'h00; mem['h5FBB]=8'h00;
    mem['h5FBC]=8'h00; mem['h5FBD]=8'h00; mem['h5FBE]=8'h00; mem['h5FBF]=8'h00;
    mem['h5FC0]=8'h00; mem['h5FC1]=8'h00; mem['h5FC2]=8'h00; mem['h5FC3]=8'h00;
    mem['h5FC4]=8'h00; mem['h5FC5]=8'h00; mem['h5FC6]=8'h00; mem['h5FC7]=8'h00;
    mem['h5FC8]=8'h00; mem['h5FC9]=8'h00; mem['h5FCA]=8'h00; mem['h5FCB]=8'h00;
    mem['h5FCC]=8'h00; mem['h5FCD]=8'h00; mem['h5FCE]=8'h00; mem['h5FCF]=8'h00;
    mem['h5FD0]=8'h00; mem['h5FD1]=8'h00; mem['h5FD2]=8'h00; mem['h5FD3]=8'h00;
    mem['h5FD4]=8'h00; mem['h5FD5]=8'h00; mem['h5FD6]=8'h00; mem['h5FD7]=8'h00;
    mem['h5FD8]=8'h00; mem['h5FD9]=8'h00; mem['h5FDA]=8'h00; mem['h5FDB]=8'h00;
    mem['h5FDC]=8'h00; mem['h5FDD]=8'h00; mem['h5FDE]=8'h00; mem['h5FDF]=8'h00;
    mem['h5FE0]=8'h00; mem['h5FE1]=8'h00; mem['h5FE2]=8'h00; mem['h5FE3]=8'h00;
    mem['h5FE4]=8'h00; mem['h5FE5]=8'h00; mem['h5FE6]=8'h00; mem['h5FE7]=8'h00;
    mem['h5FE8]=8'h00; mem['h5FE9]=8'h00; mem['h5FEA]=8'h00; mem['h5FEB]=8'h00;
    mem['h5FEC]=8'h00; mem['h5FED]=8'h00; mem['h5FEE]=8'h00; mem['h5FEF]=8'h00;
    mem['h5FF0]=8'h00; mem['h5FF1]=8'h00; mem['h5FF2]=8'h00; mem['h5FF3]=8'h00;
    mem['h5FF4]=8'h00; mem['h5FF5]=8'h00; mem['h5FF6]=8'h00; mem['h5FF7]=8'h00;
    mem['h5FF8]=8'h00; mem['h5FF9]=8'h00; mem['h5FFA]=8'h00; mem['h5FFB]=8'h00;
    mem['h5FFC]=8'h00; mem['h5FFD]=8'h00; mem['h5FFE]=8'h00; mem['h5FFF]=8'h00;
    mem['h6000]=8'h00; mem['h6001]=8'h00; mem['h6002]=8'h00; mem['h6003]=8'h00;
    mem['h6004]=8'h00; mem['h6005]=8'h00; mem['h6006]=8'h00; mem['h6007]=8'h00;
    mem['h6008]=8'h00; mem['h6009]=8'h00; mem['h600A]=8'h00; mem['h600B]=8'h00;
    mem['h600C]=8'h00; mem['h600D]=8'h00; mem['h600E]=8'h00; mem['h600F]=8'h00;
    mem['h6010]=8'h00; mem['h6011]=8'h00; mem['h6012]=8'h00; mem['h6013]=8'h00;
    mem['h6014]=8'h00; mem['h6015]=8'h00; mem['h6016]=8'h00; mem['h6017]=8'h00;
    mem['h6018]=8'h00; mem['h6019]=8'h00; mem['h601A]=8'h00; mem['h601B]=8'h00;
    mem['h601C]=8'h00; mem['h601D]=8'h00; mem['h601E]=8'h00; mem['h601F]=8'h00;
    mem['h6020]=8'h00; mem['h6021]=8'h00; mem['h6022]=8'h00; mem['h6023]=8'h00;
    mem['h6024]=8'h00; mem['h6025]=8'h00; mem['h6026]=8'h00; mem['h6027]=8'h00;
    mem['h6028]=8'h00; mem['h6029]=8'h00; mem['h602A]=8'h00; mem['h602B]=8'h00;
    mem['h602C]=8'h00; mem['h602D]=8'h00; mem['h602E]=8'h00; mem['h602F]=8'h00;
    mem['h6030]=8'h00; mem['h6031]=8'h00; mem['h6032]=8'h00; mem['h6033]=8'h00;
    mem['h6034]=8'h00; mem['h6035]=8'h00; mem['h6036]=8'h00; mem['h6037]=8'h00;
    mem['h6038]=8'h00; mem['h6039]=8'h00; mem['h603A]=8'h00; mem['h603B]=8'h00;
    mem['h603C]=8'h00; mem['h603D]=8'h00; mem['h603E]=8'h00; mem['h603F]=8'h00;
    mem['h6040]=8'h00; mem['h6041]=8'h00; mem['h6042]=8'h00; mem['h6043]=8'h00;
    mem['h6044]=8'h00; mem['h6045]=8'h00; mem['h6046]=8'h00; mem['h6047]=8'h00;
    mem['h6048]=8'h00; mem['h6049]=8'h00; mem['h604A]=8'h00; mem['h604B]=8'h00;
    mem['h604C]=8'h00; mem['h604D]=8'h00; mem['h604E]=8'h00; mem['h604F]=8'h00;
    mem['h6050]=8'h00; mem['h6051]=8'h00; mem['h6052]=8'h00; mem['h6053]=8'h00;
    mem['h6054]=8'h00; mem['h6055]=8'h00; mem['h6056]=8'h00; mem['h6057]=8'h00;
    mem['h6058]=8'h00; mem['h6059]=8'h00; mem['h605A]=8'h00; mem['h605B]=8'h00;
    mem['h605C]=8'h00; mem['h605D]=8'h00; mem['h605E]=8'h00; mem['h605F]=8'h00;
    mem['h6060]=8'h00; mem['h6061]=8'h00; mem['h6062]=8'h00; mem['h6063]=8'h00;
    mem['h6064]=8'h00; mem['h6065]=8'h00; mem['h6066]=8'h00; mem['h6067]=8'h00;
    mem['h6068]=8'h00; mem['h6069]=8'h00; mem['h606A]=8'h00; mem['h606B]=8'h00;
    mem['h606C]=8'h00; mem['h606D]=8'h00; mem['h606E]=8'h00; mem['h606F]=8'h00;
    mem['h6070]=8'h00; mem['h6071]=8'h00; mem['h6072]=8'h00; mem['h6073]=8'h00;
    mem['h6074]=8'h00; mem['h6075]=8'h00; mem['h6076]=8'h00; mem['h6077]=8'h00;
    mem['h6078]=8'h00; mem['h6079]=8'h00; mem['h607A]=8'h00; mem['h607B]=8'h00;
    mem['h607C]=8'h00; mem['h607D]=8'h00; mem['h607E]=8'h00; mem['h607F]=8'h00;
    mem['h6080]=8'h00; mem['h6081]=8'h00; mem['h6082]=8'h00; mem['h6083]=8'h00;
    mem['h6084]=8'h00; mem['h6085]=8'h00; mem['h6086]=8'h00; mem['h6087]=8'h00;
    mem['h6088]=8'h00; mem['h6089]=8'h00; mem['h608A]=8'h00; mem['h608B]=8'h00;
    mem['h608C]=8'h00; mem['h608D]=8'h00; mem['h608E]=8'h00; mem['h608F]=8'h00;
    mem['h6090]=8'h00; mem['h6091]=8'h00; mem['h6092]=8'h00; mem['h6093]=8'h00;
    mem['h6094]=8'h00; mem['h6095]=8'h00; mem['h6096]=8'h00; mem['h6097]=8'h00;
    mem['h6098]=8'h00; mem['h6099]=8'h00; mem['h609A]=8'h00; mem['h609B]=8'h00;
    mem['h609C]=8'h00; mem['h609D]=8'h00; mem['h609E]=8'h00; mem['h609F]=8'h00;
    mem['h60A0]=8'h00; mem['h60A1]=8'h00; mem['h60A2]=8'h00; mem['h60A3]=8'h00;
    mem['h60A4]=8'h00; mem['h60A5]=8'h00; mem['h60A6]=8'h00; mem['h60A7]=8'h00;
    mem['h60A8]=8'h00; mem['h60A9]=8'h00; mem['h60AA]=8'h00; mem['h60AB]=8'h00;
    mem['h60AC]=8'h00; mem['h60AD]=8'h00; mem['h60AE]=8'h00; mem['h60AF]=8'h00;
    mem['h60B0]=8'h00; mem['h60B1]=8'h00; mem['h60B2]=8'h00; mem['h60B3]=8'h00;
    mem['h60B4]=8'h00; mem['h60B5]=8'h00; mem['h60B6]=8'h00; mem['h60B7]=8'h00;
    mem['h60B8]=8'h00; mem['h60B9]=8'h00; mem['h60BA]=8'h00; mem['h60BB]=8'h00;
    mem['h60BC]=8'h00; mem['h60BD]=8'h00; mem['h60BE]=8'h00; mem['h60BF]=8'h00;
    mem['h60C0]=8'h00; mem['h60C1]=8'h00; mem['h60C2]=8'h00; mem['h60C3]=8'h00;
    mem['h60C4]=8'h00; mem['h60C5]=8'h00; mem['h60C6]=8'h00; mem['h60C7]=8'h00;
    mem['h60C8]=8'h00; mem['h60C9]=8'h00; mem['h60CA]=8'h00; mem['h60CB]=8'h00;
    mem['h60CC]=8'h00; mem['h60CD]=8'h00; mem['h60CE]=8'h00; mem['h60CF]=8'h00;
    mem['h60D0]=8'h00; mem['h60D1]=8'h00; mem['h60D2]=8'h00; mem['h60D3]=8'h00;
    mem['h60D4]=8'h00; mem['h60D5]=8'h00; mem['h60D6]=8'h00; mem['h60D7]=8'h00;
    mem['h60D8]=8'h00; mem['h60D9]=8'h00; mem['h60DA]=8'h00; mem['h60DB]=8'h00;
    mem['h60DC]=8'h00; mem['h60DD]=8'h00; mem['h60DE]=8'h00; mem['h60DF]=8'h00;
    mem['h60E0]=8'h00; mem['h60E1]=8'h00; mem['h60E2]=8'h00; mem['h60E3]=8'h00;
    mem['h60E4]=8'h00; mem['h60E5]=8'h00; mem['h60E6]=8'h00; mem['h60E7]=8'h00;
    mem['h60E8]=8'h00; mem['h60E9]=8'h00; mem['h60EA]=8'h00; mem['h60EB]=8'h00;
    mem['h60EC]=8'h00; mem['h60ED]=8'h00; mem['h60EE]=8'h00; mem['h60EF]=8'h00;
    mem['h60F0]=8'h00; mem['h60F1]=8'h00; mem['h60F2]=8'h00; mem['h60F3]=8'h00;
    mem['h60F4]=8'h00; mem['h60F5]=8'h00; mem['h60F6]=8'h00; mem['h60F7]=8'h00;
    mem['h60F8]=8'h00; mem['h60F9]=8'h00; mem['h60FA]=8'h00; mem['h60FB]=8'h00;
    mem['h60FC]=8'h00; mem['h60FD]=8'h00; mem['h60FE]=8'h00; mem['h60FF]=8'h00;
    mem['h6100]=8'h00; mem['h6101]=8'h00; mem['h6102]=8'h00; mem['h6103]=8'h00;
    mem['h6104]=8'h00; mem['h6105]=8'h00; mem['h6106]=8'h00; mem['h6107]=8'h00;
    mem['h6108]=8'h00; mem['h6109]=8'h00; mem['h610A]=8'h00; mem['h610B]=8'h00;
    mem['h610C]=8'h00; mem['h610D]=8'h00; mem['h610E]=8'h00; mem['h610F]=8'h00;
    mem['h6110]=8'h00; mem['h6111]=8'h00; mem['h6112]=8'h00; mem['h6113]=8'h00;
    mem['h6114]=8'h00; mem['h6115]=8'h00; mem['h6116]=8'h00; mem['h6117]=8'h00;
    mem['h6118]=8'h00; mem['h6119]=8'h00; mem['h611A]=8'h00; mem['h611B]=8'h00;
    mem['h611C]=8'h00; mem['h611D]=8'h00; mem['h611E]=8'h00; mem['h611F]=8'h00;
    mem['h6120]=8'h00; mem['h6121]=8'h00; mem['h6122]=8'h00; mem['h6123]=8'h00;
    mem['h6124]=8'h00; mem['h6125]=8'h00; mem['h6126]=8'h00; mem['h6127]=8'h00;
    mem['h6128]=8'h00; mem['h6129]=8'h00; mem['h612A]=8'h00; mem['h612B]=8'h00;
    mem['h612C]=8'h00; mem['h612D]=8'h00; mem['h612E]=8'h00; mem['h612F]=8'h00;
    mem['h6130]=8'h00; mem['h6131]=8'h00; mem['h6132]=8'h00; mem['h6133]=8'h00;
    mem['h6134]=8'h00; mem['h6135]=8'h00; mem['h6136]=8'h00; mem['h6137]=8'h00;
    mem['h6138]=8'h00; mem['h6139]=8'h00; mem['h613A]=8'h00; mem['h613B]=8'h00;
    mem['h613C]=8'h00; mem['h613D]=8'h00; mem['h613E]=8'h00; mem['h613F]=8'h00;
    mem['h6140]=8'h00; mem['h6141]=8'h00; mem['h6142]=8'h00; mem['h6143]=8'h00;
    mem['h6144]=8'h00; mem['h6145]=8'h00; mem['h6146]=8'h00; mem['h6147]=8'h00;
    mem['h6148]=8'h00; mem['h6149]=8'h00; mem['h614A]=8'h00; mem['h614B]=8'h00;
    mem['h614C]=8'h00; mem['h614D]=8'h00; mem['h614E]=8'h00; mem['h614F]=8'h00;
    mem['h6150]=8'h00; mem['h6151]=8'h00; mem['h6152]=8'h00; mem['h6153]=8'h00;
    mem['h6154]=8'h00; mem['h6155]=8'h00; mem['h6156]=8'h00; mem['h6157]=8'h00;
    mem['h6158]=8'h00; mem['h6159]=8'h00; mem['h615A]=8'h00; mem['h615B]=8'h00;
    mem['h615C]=8'h00; mem['h615D]=8'h00; mem['h615E]=8'h00; mem['h615F]=8'h00;
    mem['h6160]=8'h00; mem['h6161]=8'h00; mem['h6162]=8'h00; mem['h6163]=8'h00;
    mem['h6164]=8'h00; mem['h6165]=8'h00; mem['h6166]=8'h00; mem['h6167]=8'h00;
    mem['h6168]=8'h00; mem['h6169]=8'h00; mem['h616A]=8'h00; mem['h616B]=8'h00;
    mem['h616C]=8'h00; mem['h616D]=8'h00; mem['h616E]=8'h00; mem['h616F]=8'h00;
    mem['h6170]=8'h00; mem['h6171]=8'h00; mem['h6172]=8'h00; mem['h6173]=8'h00;
    mem['h6174]=8'h00; mem['h6175]=8'h00; mem['h6176]=8'h00; mem['h6177]=8'h00;
    mem['h6178]=8'h00; mem['h6179]=8'h00; mem['h617A]=8'h00; mem['h617B]=8'h00;
    mem['h617C]=8'h00; mem['h617D]=8'h00; mem['h617E]=8'h00; mem['h617F]=8'h00;
    mem['h6180]=8'h00; mem['h6181]=8'h00; mem['h6182]=8'h00; mem['h6183]=8'h00;
    mem['h6184]=8'h00; mem['h6185]=8'h00; mem['h6186]=8'h00; mem['h6187]=8'h00;
    mem['h6188]=8'h00; mem['h6189]=8'h00; mem['h618A]=8'h00; mem['h618B]=8'h00;
    mem['h618C]=8'h00; mem['h618D]=8'h00; mem['h618E]=8'h00; mem['h618F]=8'h00;
    mem['h6190]=8'h00; mem['h6191]=8'h00; mem['h6192]=8'h00; mem['h6193]=8'h00;
    mem['h6194]=8'h00; mem['h6195]=8'h00; mem['h6196]=8'h00; mem['h6197]=8'h00;
    mem['h6198]=8'h00; mem['h6199]=8'h00; mem['h619A]=8'h00; mem['h619B]=8'h00;
    mem['h619C]=8'h00; mem['h619D]=8'h00; mem['h619E]=8'h00; mem['h619F]=8'h00;
    mem['h61A0]=8'h00; mem['h61A1]=8'h00; mem['h61A2]=8'h00; mem['h61A3]=8'h00;
    mem['h61A4]=8'h00; mem['h61A5]=8'h00; mem['h61A6]=8'h00; mem['h61A7]=8'h00;
    mem['h61A8]=8'h00; mem['h61A9]=8'h00; mem['h61AA]=8'h00; mem['h61AB]=8'h00;
    mem['h61AC]=8'h00; mem['h61AD]=8'h00; mem['h61AE]=8'h00; mem['h61AF]=8'h00;
    mem['h61B0]=8'h00; mem['h61B1]=8'h00; mem['h61B2]=8'h00; mem['h61B3]=8'h00;
    mem['h61B4]=8'h00; mem['h61B5]=8'h00; mem['h61B6]=8'h00; mem['h61B7]=8'h00;
    mem['h61B8]=8'h00; mem['h61B9]=8'h00; mem['h61BA]=8'h00; mem['h61BB]=8'h00;
    mem['h61BC]=8'h00; mem['h61BD]=8'h00; mem['h61BE]=8'h00; mem['h61BF]=8'h00;
    mem['h61C0]=8'h00; mem['h61C1]=8'h00; mem['h61C2]=8'h00; mem['h61C3]=8'h00;
    mem['h61C4]=8'h00; mem['h61C5]=8'h00; mem['h61C6]=8'h00; mem['h61C7]=8'h00;
    mem['h61C8]=8'h00; mem['h61C9]=8'h00; mem['h61CA]=8'h00; mem['h61CB]=8'h00;
    mem['h61CC]=8'h00; mem['h61CD]=8'h00; mem['h61CE]=8'h00; mem['h61CF]=8'h00;
    mem['h61D0]=8'h00; mem['h61D1]=8'h00; mem['h61D2]=8'h00; mem['h61D3]=8'h00;
    mem['h61D4]=8'h00; mem['h61D5]=8'h00; mem['h61D6]=8'h00; mem['h61D7]=8'h00;
    mem['h61D8]=8'h00; mem['h61D9]=8'h00; mem['h61DA]=8'h00; mem['h61DB]=8'h00;
    mem['h61DC]=8'h00; mem['h61DD]=8'h00; mem['h61DE]=8'h00; mem['h61DF]=8'h00;
    mem['h61E0]=8'h00; mem['h61E1]=8'h00; mem['h61E2]=8'h00; mem['h61E3]=8'h00;
    mem['h61E4]=8'h00; mem['h61E5]=8'h00; mem['h61E6]=8'h00; mem['h61E7]=8'h00;
    mem['h61E8]=8'h00; mem['h61E9]=8'h00; mem['h61EA]=8'h00; mem['h61EB]=8'h00;
    mem['h61EC]=8'h00; mem['h61ED]=8'h00; mem['h61EE]=8'h00; mem['h61EF]=8'h00;
    mem['h61F0]=8'h00; mem['h61F1]=8'h00; mem['h61F2]=8'h00; mem['h61F3]=8'h00;
    mem['h61F4]=8'h00; mem['h61F5]=8'h00; mem['h61F6]=8'h00; mem['h61F7]=8'h00;
    mem['h61F8]=8'h00; mem['h61F9]=8'h00; mem['h61FA]=8'h00; mem['h61FB]=8'h00;
    mem['h61FC]=8'h00; mem['h61FD]=8'h00; mem['h61FE]=8'h00; mem['h61FF]=8'h00;
    mem['h6200]=8'h00; mem['h6201]=8'h00; mem['h6202]=8'h00; mem['h6203]=8'h00;
    mem['h6204]=8'h00; mem['h6205]=8'h00; mem['h6206]=8'h00; mem['h6207]=8'h00;
    mem['h6208]=8'h00; mem['h6209]=8'h00; mem['h620A]=8'h00; mem['h620B]=8'h00;
    mem['h620C]=8'h00; mem['h620D]=8'h00; mem['h620E]=8'h00; mem['h620F]=8'h00;
    mem['h6210]=8'h00; mem['h6211]=8'h00; mem['h6212]=8'h00; mem['h6213]=8'h00;
    mem['h6214]=8'h00; mem['h6215]=8'h00; mem['h6216]=8'h00; mem['h6217]=8'h00;
    mem['h6218]=8'h00; mem['h6219]=8'h00; mem['h621A]=8'h00; mem['h621B]=8'h00;
    mem['h621C]=8'h00; mem['h621D]=8'h00; mem['h621E]=8'h00; mem['h621F]=8'h00;
    mem['h6220]=8'h00; mem['h6221]=8'h00; mem['h6222]=8'h00; mem['h6223]=8'h00;
    mem['h6224]=8'h00; mem['h6225]=8'h00; mem['h6226]=8'h00; mem['h6227]=8'h00;
    mem['h6228]=8'h00; mem['h6229]=8'h00; mem['h622A]=8'h00; mem['h622B]=8'h00;
    mem['h622C]=8'h00; mem['h622D]=8'h00; mem['h622E]=8'h00; mem['h622F]=8'h00;
    mem['h6230]=8'h00; mem['h6231]=8'h00; mem['h6232]=8'h00; mem['h6233]=8'h00;
    mem['h6234]=8'h00; mem['h6235]=8'h00; mem['h6236]=8'h00; mem['h6237]=8'h00;
    mem['h6238]=8'h00; mem['h6239]=8'h00; mem['h623A]=8'h00; mem['h623B]=8'h00;
    mem['h623C]=8'h00; mem['h623D]=8'h00; mem['h623E]=8'h00; mem['h623F]=8'h00;
    mem['h6240]=8'h00; mem['h6241]=8'h00; mem['h6242]=8'h00; mem['h6243]=8'h00;
    mem['h6244]=8'h00; mem['h6245]=8'h00; mem['h6246]=8'h00; mem['h6247]=8'h00;
    mem['h6248]=8'h00; mem['h6249]=8'h00; mem['h624A]=8'h00; mem['h624B]=8'h00;
    mem['h624C]=8'h00; mem['h624D]=8'h00; mem['h624E]=8'h00; mem['h624F]=8'h00;
    mem['h6250]=8'h00; mem['h6251]=8'h00; mem['h6252]=8'h00; mem['h6253]=8'h00;
    mem['h6254]=8'h00; mem['h6255]=8'h00; mem['h6256]=8'h00; mem['h6257]=8'h00;
    mem['h6258]=8'h00; mem['h6259]=8'h00; mem['h625A]=8'h00; mem['h625B]=8'h00;
    mem['h625C]=8'h00; mem['h625D]=8'h00; mem['h625E]=8'h00; mem['h625F]=8'h00;
    mem['h6260]=8'h00; mem['h6261]=8'h00; mem['h6262]=8'h00; mem['h6263]=8'h00;
    mem['h6264]=8'h00; mem['h6265]=8'h00; mem['h6266]=8'h00; mem['h6267]=8'h00;
    mem['h6268]=8'h00; mem['h6269]=8'h00; mem['h626A]=8'h00; mem['h626B]=8'h00;
    mem['h626C]=8'h00; mem['h626D]=8'h00; mem['h626E]=8'h00; mem['h626F]=8'h00;
    mem['h6270]=8'h00; mem['h6271]=8'h00; mem['h6272]=8'h00; mem['h6273]=8'h00;
    mem['h6274]=8'h00; mem['h6275]=8'h00; mem['h6276]=8'h00; mem['h6277]=8'h00;
    mem['h6278]=8'h00; mem['h6279]=8'h00; mem['h627A]=8'h00; mem['h627B]=8'h00;
    mem['h627C]=8'h00; mem['h627D]=8'h00; mem['h627E]=8'h00; mem['h627F]=8'h00;
    mem['h6280]=8'h00; mem['h6281]=8'h00; mem['h6282]=8'h00; mem['h6283]=8'h00;
    mem['h6284]=8'h00; mem['h6285]=8'h00; mem['h6286]=8'h00; mem['h6287]=8'h00;
    mem['h6288]=8'h00; mem['h6289]=8'h00; mem['h628A]=8'h00; mem['h628B]=8'h00;
    mem['h628C]=8'h00; mem['h628D]=8'h00; mem['h628E]=8'h00; mem['h628F]=8'h00;
    mem['h6290]=8'h00; mem['h6291]=8'h00; mem['h6292]=8'h00; mem['h6293]=8'h00;
    mem['h6294]=8'h00; mem['h6295]=8'h00; mem['h6296]=8'h00; mem['h6297]=8'h00;
    mem['h6298]=8'h00; mem['h6299]=8'h00; mem['h629A]=8'h00; mem['h629B]=8'h00;
    mem['h629C]=8'h00; mem['h629D]=8'h00; mem['h629E]=8'h00; mem['h629F]=8'h00;
    mem['h62A0]=8'h00; mem['h62A1]=8'h00; mem['h62A2]=8'h00; mem['h62A3]=8'h00;
    mem['h62A4]=8'h00; mem['h62A5]=8'h00; mem['h62A6]=8'h00; mem['h62A7]=8'h00;
    mem['h62A8]=8'h00; mem['h62A9]=8'h00; mem['h62AA]=8'h00; mem['h62AB]=8'h00;
    mem['h62AC]=8'h00; mem['h62AD]=8'h00; mem['h62AE]=8'h00; mem['h62AF]=8'h00;
    mem['h62B0]=8'h00; mem['h62B1]=8'h00; mem['h62B2]=8'h00; mem['h62B3]=8'h00;
    mem['h62B4]=8'h00; mem['h62B5]=8'h00; mem['h62B6]=8'h00; mem['h62B7]=8'h00;
    mem['h62B8]=8'h00; mem['h62B9]=8'h00; mem['h62BA]=8'h00; mem['h62BB]=8'h00;
    mem['h62BC]=8'h00; mem['h62BD]=8'h00; mem['h62BE]=8'h00; mem['h62BF]=8'h00;
    mem['h62C0]=8'h00; mem['h62C1]=8'h00; mem['h62C2]=8'h00; mem['h62C3]=8'h00;
    mem['h62C4]=8'h00; mem['h62C5]=8'h00; mem['h62C6]=8'h00; mem['h62C7]=8'h00;
    mem['h62C8]=8'h00; mem['h62C9]=8'h00; mem['h62CA]=8'h00; mem['h62CB]=8'h00;
    mem['h62CC]=8'h00; mem['h62CD]=8'h00; mem['h62CE]=8'h00; mem['h62CF]=8'h00;
    mem['h62D0]=8'h00; mem['h62D1]=8'h00; mem['h62D2]=8'h00; mem['h62D3]=8'h00;
    mem['h62D4]=8'h00; mem['h62D5]=8'h00; mem['h62D6]=8'h00; mem['h62D7]=8'h00;
    mem['h62D8]=8'h00; mem['h62D9]=8'h00; mem['h62DA]=8'h00; mem['h62DB]=8'h00;
    mem['h62DC]=8'h00; mem['h62DD]=8'h00; mem['h62DE]=8'h00; mem['h62DF]=8'h00;
    mem['h62E0]=8'h00; mem['h62E1]=8'h00; mem['h62E2]=8'h00; mem['h62E3]=8'h00;
    mem['h62E4]=8'h00; mem['h62E5]=8'h00; mem['h62E6]=8'h00; mem['h62E7]=8'h00;
    mem['h62E8]=8'h00; mem['h62E9]=8'h00; mem['h62EA]=8'h00; mem['h62EB]=8'h00;
    mem['h62EC]=8'h00; mem['h62ED]=8'h00; mem['h62EE]=8'h00; mem['h62EF]=8'h00;
    mem['h62F0]=8'h00; mem['h62F1]=8'h00; mem['h62F2]=8'h00; mem['h62F3]=8'h00;
    mem['h62F4]=8'h00; mem['h62F5]=8'h00; mem['h62F6]=8'h00; mem['h62F7]=8'h00;
    mem['h62F8]=8'h00; mem['h62F9]=8'h00; mem['h62FA]=8'h00; mem['h62FB]=8'h00;
    mem['h62FC]=8'h00; mem['h62FD]=8'h00; mem['h62FE]=8'h00; mem['h62FF]=8'h00;
    mem['h6300]=8'h00; mem['h6301]=8'h00; mem['h6302]=8'h00; mem['h6303]=8'h00;
    mem['h6304]=8'h00; mem['h6305]=8'h00; mem['h6306]=8'h00; mem['h6307]=8'h00;
    mem['h6308]=8'h00; mem['h6309]=8'h00; mem['h630A]=8'h00; mem['h630B]=8'h00;
    mem['h630C]=8'h00; mem['h630D]=8'h00; mem['h630E]=8'h00; mem['h630F]=8'h00;
    mem['h6310]=8'h00; mem['h6311]=8'h00; mem['h6312]=8'h00; mem['h6313]=8'h00;
    mem['h6314]=8'h00; mem['h6315]=8'h00; mem['h6316]=8'h00; mem['h6317]=8'h00;
    mem['h6318]=8'h00; mem['h6319]=8'h00; mem['h631A]=8'h00; mem['h631B]=8'h00;
    mem['h631C]=8'h00; mem['h631D]=8'h00; mem['h631E]=8'h00; mem['h631F]=8'h00;
    mem['h6320]=8'h00; mem['h6321]=8'h00; mem['h6322]=8'h00; mem['h6323]=8'h00;
    mem['h6324]=8'h00; mem['h6325]=8'h00; mem['h6326]=8'h00; mem['h6327]=8'h00;
    mem['h6328]=8'h00; mem['h6329]=8'h00; mem['h632A]=8'h00; mem['h632B]=8'h00;
    mem['h632C]=8'h00; mem['h632D]=8'h00; mem['h632E]=8'h00; mem['h632F]=8'h00;
    mem['h6330]=8'h00; mem['h6331]=8'h00; mem['h6332]=8'h00; mem['h6333]=8'h00;
    mem['h6334]=8'h00; mem['h6335]=8'h00; mem['h6336]=8'h00; mem['h6337]=8'h00;
    mem['h6338]=8'h00; mem['h6339]=8'h00; mem['h633A]=8'h00; mem['h633B]=8'h00;
    mem['h633C]=8'h00; mem['h633D]=8'h00; mem['h633E]=8'h00; mem['h633F]=8'h00;
    mem['h6340]=8'h00; mem['h6341]=8'h00; mem['h6342]=8'h00; mem['h6343]=8'h00;
    mem['h6344]=8'h00; mem['h6345]=8'h00; mem['h6346]=8'h00; mem['h6347]=8'h00;
    mem['h6348]=8'h00; mem['h6349]=8'h00; mem['h634A]=8'h00; mem['h634B]=8'h00;
    mem['h634C]=8'h00; mem['h634D]=8'h00; mem['h634E]=8'h00; mem['h634F]=8'h00;
    mem['h6350]=8'h00; mem['h6351]=8'h00; mem['h6352]=8'h00; mem['h6353]=8'h00;
    mem['h6354]=8'h00; mem['h6355]=8'h00; mem['h6356]=8'h00; mem['h6357]=8'h00;
    mem['h6358]=8'h00; mem['h6359]=8'h00; mem['h635A]=8'h00; mem['h635B]=8'h00;
    mem['h635C]=8'h00; mem['h635D]=8'h00; mem['h635E]=8'h00; mem['h635F]=8'h00;
    mem['h6360]=8'h00; mem['h6361]=8'h00; mem['h6362]=8'h00; mem['h6363]=8'h00;
    mem['h6364]=8'h00; mem['h6365]=8'h00; mem['h6366]=8'h00; mem['h6367]=8'h00;
    mem['h6368]=8'h00; mem['h6369]=8'h00; mem['h636A]=8'h00; mem['h636B]=8'h00;
    mem['h636C]=8'h00; mem['h636D]=8'h00; mem['h636E]=8'h00; mem['h636F]=8'h00;
    mem['h6370]=8'h00; mem['h6371]=8'h00; mem['h6372]=8'h00; mem['h6373]=8'h00;
    mem['h6374]=8'h00; mem['h6375]=8'h00; mem['h6376]=8'h00; mem['h6377]=8'h00;
    mem['h6378]=8'h00; mem['h6379]=8'h00; mem['h637A]=8'h00; mem['h637B]=8'h00;
    mem['h637C]=8'h00; mem['h637D]=8'h00; mem['h637E]=8'h00; mem['h637F]=8'h00;
    mem['h6380]=8'h00; mem['h6381]=8'h00; mem['h6382]=8'h00; mem['h6383]=8'h00;
    mem['h6384]=8'h00; mem['h6385]=8'h00; mem['h6386]=8'h00; mem['h6387]=8'h00;
    mem['h6388]=8'h00; mem['h6389]=8'h00; mem['h638A]=8'h00; mem['h638B]=8'h00;
    mem['h638C]=8'h00; mem['h638D]=8'h00; mem['h638E]=8'h00; mem['h638F]=8'h00;
    mem['h6390]=8'h00; mem['h6391]=8'h00; mem['h6392]=8'h00; mem['h6393]=8'h00;
    mem['h6394]=8'h00; mem['h6395]=8'h00; mem['h6396]=8'h00; mem['h6397]=8'h00;
    mem['h6398]=8'h00; mem['h6399]=8'h00; mem['h639A]=8'h00; mem['h639B]=8'h00;
    mem['h639C]=8'h00; mem['h639D]=8'h00; mem['h639E]=8'h00; mem['h639F]=8'h00;
    mem['h63A0]=8'h00; mem['h63A1]=8'h00; mem['h63A2]=8'h00; mem['h63A3]=8'h00;
    mem['h63A4]=8'h00; mem['h63A5]=8'h00; mem['h63A6]=8'h00; mem['h63A7]=8'h00;
    mem['h63A8]=8'h00; mem['h63A9]=8'h00; mem['h63AA]=8'h00; mem['h63AB]=8'h00;
    mem['h63AC]=8'h00; mem['h63AD]=8'h00; mem['h63AE]=8'h00; mem['h63AF]=8'h00;
    mem['h63B0]=8'h00; mem['h63B1]=8'h00; mem['h63B2]=8'h00; mem['h63B3]=8'h00;
    mem['h63B4]=8'h00; mem['h63B5]=8'h00; mem['h63B6]=8'h00; mem['h63B7]=8'h00;
    mem['h63B8]=8'h00; mem['h63B9]=8'h00; mem['h63BA]=8'h00; mem['h63BB]=8'h00;
    mem['h63BC]=8'h00; mem['h63BD]=8'h00; mem['h63BE]=8'h00; mem['h63BF]=8'h00;
    mem['h63C0]=8'h00; mem['h63C1]=8'h00; mem['h63C2]=8'h00; mem['h63C3]=8'h00;
    mem['h63C4]=8'h00; mem['h63C5]=8'h00; mem['h63C6]=8'h00; mem['h63C7]=8'h00;
    mem['h63C8]=8'h00; mem['h63C9]=8'h00; mem['h63CA]=8'h00; mem['h63CB]=8'h00;
    mem['h63CC]=8'h00; mem['h63CD]=8'h00; mem['h63CE]=8'h00; mem['h63CF]=8'h00;
    mem['h63D0]=8'h00; mem['h63D1]=8'h00; mem['h63D2]=8'h00; mem['h63D3]=8'h00;
    mem['h63D4]=8'h00; mem['h63D5]=8'h00; mem['h63D6]=8'h00; mem['h63D7]=8'h00;
    mem['h63D8]=8'h00; mem['h63D9]=8'h00; mem['h63DA]=8'h00; mem['h63DB]=8'h00;
    mem['h63DC]=8'h00; mem['h63DD]=8'h00; mem['h63DE]=8'h00; mem['h63DF]=8'h00;
    mem['h63E0]=8'h00; mem['h63E1]=8'h00; mem['h63E2]=8'h00; mem['h63E3]=8'h00;
    mem['h63E4]=8'h00; mem['h63E5]=8'h00; mem['h63E6]=8'h00; mem['h63E7]=8'h00;
    mem['h63E8]=8'h00; mem['h63E9]=8'h00; mem['h63EA]=8'h00; mem['h63EB]=8'h00;
    mem['h63EC]=8'h00; mem['h63ED]=8'h00; mem['h63EE]=8'h00; mem['h63EF]=8'h00;
    mem['h63F0]=8'h00; mem['h63F1]=8'h00; mem['h63F2]=8'h00; mem['h63F3]=8'h00;
    mem['h63F4]=8'h00; mem['h63F5]=8'h00; mem['h63F6]=8'h00; mem['h63F7]=8'h00;
    mem['h63F8]=8'h00; mem['h63F9]=8'h00; mem['h63FA]=8'h00; mem['h63FB]=8'h00;
    mem['h63FC]=8'h00; mem['h63FD]=8'h00; mem['h63FE]=8'h00; mem['h63FF]=8'h00;
    mem['h6400]=8'h00; mem['h6401]=8'h00; mem['h6402]=8'h00; mem['h6403]=8'h00;
    mem['h6404]=8'h00; mem['h6405]=8'h00; mem['h6406]=8'h00; mem['h6407]=8'h00;
    mem['h6408]=8'h00; mem['h6409]=8'h00; mem['h640A]=8'h00; mem['h640B]=8'h00;
    mem['h640C]=8'h00; mem['h640D]=8'h00; mem['h640E]=8'h00; mem['h640F]=8'h00;
    mem['h6410]=8'h00; mem['h6411]=8'h00; mem['h6412]=8'h00; mem['h6413]=8'h00;
    mem['h6414]=8'h00; mem['h6415]=8'h00; mem['h6416]=8'h00; mem['h6417]=8'h00;
    mem['h6418]=8'h00; mem['h6419]=8'h00; mem['h641A]=8'h00; mem['h641B]=8'h00;
    mem['h641C]=8'h00; mem['h641D]=8'h00; mem['h641E]=8'h00; mem['h641F]=8'h00;
    mem['h6420]=8'h00; mem['h6421]=8'h00; mem['h6422]=8'h00; mem['h6423]=8'h00;
    mem['h6424]=8'h00; mem['h6425]=8'h00; mem['h6426]=8'h00; mem['h6427]=8'h00;
    mem['h6428]=8'h00; mem['h6429]=8'h00; mem['h642A]=8'h00; mem['h642B]=8'h00;
    mem['h642C]=8'h00; mem['h642D]=8'h00; mem['h642E]=8'h00; mem['h642F]=8'h00;
    mem['h6430]=8'h00; mem['h6431]=8'h00; mem['h6432]=8'h00; mem['h6433]=8'h00;
    mem['h6434]=8'h00; mem['h6435]=8'h00; mem['h6436]=8'h00; mem['h6437]=8'h00;
    mem['h6438]=8'h00; mem['h6439]=8'h00; mem['h643A]=8'h00; mem['h643B]=8'h00;
    mem['h643C]=8'h00; mem['h643D]=8'h00; mem['h643E]=8'h00; mem['h643F]=8'h00;
    mem['h6440]=8'h00; mem['h6441]=8'h00; mem['h6442]=8'h00; mem['h6443]=8'h00;
    mem['h6444]=8'h00; mem['h6445]=8'h00; mem['h6446]=8'h00; mem['h6447]=8'h00;
    mem['h6448]=8'h00; mem['h6449]=8'h00; mem['h644A]=8'h00; mem['h644B]=8'h00;
    mem['h644C]=8'h00; mem['h644D]=8'h00; mem['h644E]=8'h00; mem['h644F]=8'h00;
    mem['h6450]=8'h00; mem['h6451]=8'h00; mem['h6452]=8'h00; mem['h6453]=8'h00;
    mem['h6454]=8'h00; mem['h6455]=8'h00; mem['h6456]=8'h00; mem['h6457]=8'h00;
    mem['h6458]=8'h00; mem['h6459]=8'h00; mem['h645A]=8'h00; mem['h645B]=8'h00;
    mem['h645C]=8'h00; mem['h645D]=8'h00; mem['h645E]=8'h00; mem['h645F]=8'h00;
    mem['h6460]=8'h00; mem['h6461]=8'h00; mem['h6462]=8'h00; mem['h6463]=8'h00;
    mem['h6464]=8'h00; mem['h6465]=8'h00; mem['h6466]=8'h00; mem['h6467]=8'h00;
    mem['h6468]=8'h00; mem['h6469]=8'h00; mem['h646A]=8'h00; mem['h646B]=8'h00;
    mem['h646C]=8'h00; mem['h646D]=8'h00; mem['h646E]=8'h00; mem['h646F]=8'h00;
    mem['h6470]=8'h00; mem['h6471]=8'h00; mem['h6472]=8'h00; mem['h6473]=8'h00;
    mem['h6474]=8'h00; mem['h6475]=8'h00; mem['h6476]=8'h00; mem['h6477]=8'h00;
    mem['h6478]=8'h00; mem['h6479]=8'h00; mem['h647A]=8'h00; mem['h647B]=8'h00;
    mem['h647C]=8'h00; mem['h647D]=8'h00; mem['h647E]=8'h00; mem['h647F]=8'h00;
    mem['h6480]=8'h00; mem['h6481]=8'h00; mem['h6482]=8'h00; mem['h6483]=8'h00;
    mem['h6484]=8'h00; mem['h6485]=8'h00; mem['h6486]=8'h00; mem['h6487]=8'h00;
    mem['h6488]=8'h00; mem['h6489]=8'h00; mem['h648A]=8'h00; mem['h648B]=8'h00;
    mem['h648C]=8'h00; mem['h648D]=8'h00; mem['h648E]=8'h00; mem['h648F]=8'h00;
    mem['h6490]=8'h00; mem['h6491]=8'h00; mem['h6492]=8'h00; mem['h6493]=8'h00;
    mem['h6494]=8'h00; mem['h6495]=8'h00; mem['h6496]=8'h00; mem['h6497]=8'h00;
    mem['h6498]=8'h00; mem['h6499]=8'h00; mem['h649A]=8'h00; mem['h649B]=8'h00;
    mem['h649C]=8'h00; mem['h649D]=8'h00; mem['h649E]=8'h00; mem['h649F]=8'h00;
    mem['h64A0]=8'h00; mem['h64A1]=8'h00; mem['h64A2]=8'h00; mem['h64A3]=8'h00;
    mem['h64A4]=8'h00; mem['h64A5]=8'h00; mem['h64A6]=8'h00; mem['h64A7]=8'h00;
    mem['h64A8]=8'h00; mem['h64A9]=8'h00; mem['h64AA]=8'h00; mem['h64AB]=8'h00;
    mem['h64AC]=8'h00; mem['h64AD]=8'h00; mem['h64AE]=8'h00; mem['h64AF]=8'h00;
    mem['h64B0]=8'h00; mem['h64B1]=8'h00; mem['h64B2]=8'h00; mem['h64B3]=8'h00;
    mem['h64B4]=8'h00; mem['h64B5]=8'h00; mem['h64B6]=8'h00; mem['h64B7]=8'h00;
    mem['h64B8]=8'h00; mem['h64B9]=8'h00; mem['h64BA]=8'h00; mem['h64BB]=8'h00;
    mem['h64BC]=8'h00; mem['h64BD]=8'h00; mem['h64BE]=8'h00; mem['h64BF]=8'h00;
    mem['h64C0]=8'h00; mem['h64C1]=8'h00; mem['h64C2]=8'h00; mem['h64C3]=8'h00;
    mem['h64C4]=8'h00; mem['h64C5]=8'h00; mem['h64C6]=8'h00; mem['h64C7]=8'h00;
    mem['h64C8]=8'h00; mem['h64C9]=8'h00; mem['h64CA]=8'h00; mem['h64CB]=8'h00;
    mem['h64CC]=8'h00; mem['h64CD]=8'h00; mem['h64CE]=8'h00; mem['h64CF]=8'h00;
    mem['h64D0]=8'h00; mem['h64D1]=8'h00; mem['h64D2]=8'h00; mem['h64D3]=8'h00;
    mem['h64D4]=8'h00; mem['h64D5]=8'h00; mem['h64D6]=8'h00; mem['h64D7]=8'h00;
    mem['h64D8]=8'h00; mem['h64D9]=8'h00; mem['h64DA]=8'h00; mem['h64DB]=8'h00;
    mem['h64DC]=8'h00; mem['h64DD]=8'h00; mem['h64DE]=8'h00; mem['h64DF]=8'h00;
    mem['h64E0]=8'h00; mem['h64E1]=8'h00; mem['h64E2]=8'h00; mem['h64E3]=8'h00;
    mem['h64E4]=8'h00; mem['h64E5]=8'h00; mem['h64E6]=8'h00; mem['h64E7]=8'h00;
    mem['h64E8]=8'h00; mem['h64E9]=8'h00; mem['h64EA]=8'h00; mem['h64EB]=8'h00;
    mem['h64EC]=8'h00; mem['h64ED]=8'h00; mem['h64EE]=8'h00; mem['h64EF]=8'h00;
    mem['h64F0]=8'h00; mem['h64F1]=8'h00; mem['h64F2]=8'h00; mem['h64F3]=8'h00;
    mem['h64F4]=8'h00; mem['h64F5]=8'h00; mem['h64F6]=8'h00; mem['h64F7]=8'h00;
    mem['h64F8]=8'h00; mem['h64F9]=8'h00; mem['h64FA]=8'h00; mem['h64FB]=8'h00;
    mem['h64FC]=8'h00; mem['h64FD]=8'h00; mem['h64FE]=8'h00; mem['h64FF]=8'h00;
    mem['h6500]=8'h00; mem['h6501]=8'h00; mem['h6502]=8'h00; mem['h6503]=8'h00;
    mem['h6504]=8'h00; mem['h6505]=8'h00; mem['h6506]=8'h00; mem['h6507]=8'h00;
    mem['h6508]=8'h00; mem['h6509]=8'h00; mem['h650A]=8'h00; mem['h650B]=8'h00;
    mem['h650C]=8'h00; mem['h650D]=8'h00; mem['h650E]=8'h00; mem['h650F]=8'h00;
    mem['h6510]=8'h00; mem['h6511]=8'h00; mem['h6512]=8'h00; mem['h6513]=8'h00;
    mem['h6514]=8'h00; mem['h6515]=8'h00; mem['h6516]=8'h00; mem['h6517]=8'h00;
    mem['h6518]=8'h00; mem['h6519]=8'h00; mem['h651A]=8'h00; mem['h651B]=8'h00;
    mem['h651C]=8'h00; mem['h651D]=8'h00; mem['h651E]=8'h00; mem['h651F]=8'h00;
    mem['h6520]=8'h00; mem['h6521]=8'h00; mem['h6522]=8'h00; mem['h6523]=8'h00;
    mem['h6524]=8'h00; mem['h6525]=8'h00; mem['h6526]=8'h00; mem['h6527]=8'h00;
    mem['h6528]=8'h00; mem['h6529]=8'h00; mem['h652A]=8'h00; mem['h652B]=8'h00;
    mem['h652C]=8'h00; mem['h652D]=8'h00; mem['h652E]=8'h00; mem['h652F]=8'h00;
    mem['h6530]=8'h00; mem['h6531]=8'h00; mem['h6532]=8'h00; mem['h6533]=8'h00;
    mem['h6534]=8'h00; mem['h6535]=8'h00; mem['h6536]=8'h00; mem['h6537]=8'h00;
    mem['h6538]=8'h00; mem['h6539]=8'h00; mem['h653A]=8'h00; mem['h653B]=8'h00;
    mem['h653C]=8'h00; mem['h653D]=8'h00; mem['h653E]=8'h00; mem['h653F]=8'h00;
    mem['h6540]=8'h00; mem['h6541]=8'h00; mem['h6542]=8'h00; mem['h6543]=8'h00;
    mem['h6544]=8'h00; mem['h6545]=8'h00; mem['h6546]=8'h00; mem['h6547]=8'h00;
    mem['h6548]=8'h00; mem['h6549]=8'h00; mem['h654A]=8'h00; mem['h654B]=8'h00;
    mem['h654C]=8'h00; mem['h654D]=8'h00; mem['h654E]=8'h00; mem['h654F]=8'h00;
    mem['h6550]=8'h00; mem['h6551]=8'h00; mem['h6552]=8'h00; mem['h6553]=8'h00;
    mem['h6554]=8'h00; mem['h6555]=8'h00; mem['h6556]=8'h00; mem['h6557]=8'h00;
    mem['h6558]=8'h00; mem['h6559]=8'h00; mem['h655A]=8'h00; mem['h655B]=8'h00;
    mem['h655C]=8'h00; mem['h655D]=8'h00; mem['h655E]=8'h00; mem['h655F]=8'h00;
    mem['h6560]=8'h00; mem['h6561]=8'h00; mem['h6562]=8'h00; mem['h6563]=8'h00;
    mem['h6564]=8'h00; mem['h6565]=8'h00; mem['h6566]=8'h00; mem['h6567]=8'h00;
    mem['h6568]=8'h00; mem['h6569]=8'h00; mem['h656A]=8'h00; mem['h656B]=8'h00;
    mem['h656C]=8'h00; mem['h656D]=8'h00; mem['h656E]=8'h00; mem['h656F]=8'h00;
    mem['h6570]=8'h00; mem['h6571]=8'h00; mem['h6572]=8'h00; mem['h6573]=8'h00;
    mem['h6574]=8'h00; mem['h6575]=8'h00; mem['h6576]=8'h00; mem['h6577]=8'h00;
    mem['h6578]=8'h00; mem['h6579]=8'h00; mem['h657A]=8'h00; mem['h657B]=8'h00;
    mem['h657C]=8'h00; mem['h657D]=8'h00; mem['h657E]=8'h00; mem['h657F]=8'h00;
    mem['h6580]=8'h00; mem['h6581]=8'h00; mem['h6582]=8'h00; mem['h6583]=8'h00;
    mem['h6584]=8'h00; mem['h6585]=8'h00; mem['h6586]=8'h00; mem['h6587]=8'h00;
    mem['h6588]=8'h00; mem['h6589]=8'h00; mem['h658A]=8'h00; mem['h658B]=8'h00;
    mem['h658C]=8'h00; mem['h658D]=8'h00; mem['h658E]=8'h00; mem['h658F]=8'h00;
    mem['h6590]=8'h00; mem['h6591]=8'h00; mem['h6592]=8'h00; mem['h6593]=8'h00;
    mem['h6594]=8'h00; mem['h6595]=8'h00; mem['h6596]=8'h00; mem['h6597]=8'h00;
    mem['h6598]=8'h00; mem['h6599]=8'h00; mem['h659A]=8'h00; mem['h659B]=8'h00;
    mem['h659C]=8'h00; mem['h659D]=8'h00; mem['h659E]=8'h00; mem['h659F]=8'h00;
    mem['h65A0]=8'h00; mem['h65A1]=8'h00; mem['h65A2]=8'h00; mem['h65A3]=8'h00;
    mem['h65A4]=8'h00; mem['h65A5]=8'h00; mem['h65A6]=8'h00; mem['h65A7]=8'h00;
    mem['h65A8]=8'h00; mem['h65A9]=8'h00; mem['h65AA]=8'h00; mem['h65AB]=8'h00;
    mem['h65AC]=8'h00; mem['h65AD]=8'h00; mem['h65AE]=8'h00; mem['h65AF]=8'h00;
    mem['h65B0]=8'h00; mem['h65B1]=8'h00; mem['h65B2]=8'h00; mem['h65B3]=8'h00;
    mem['h65B4]=8'h00; mem['h65B5]=8'h00; mem['h65B6]=8'h00; mem['h65B7]=8'h00;
    mem['h65B8]=8'h00; mem['h65B9]=8'h00; mem['h65BA]=8'h00; mem['h65BB]=8'h00;
    mem['h65BC]=8'h00; mem['h65BD]=8'h00; mem['h65BE]=8'h00; mem['h65BF]=8'h00;
    mem['h65C0]=8'h00; mem['h65C1]=8'h00; mem['h65C2]=8'h00; mem['h65C3]=8'h00;
    mem['h65C4]=8'h00; mem['h65C5]=8'h00; mem['h65C6]=8'h00; mem['h65C7]=8'h00;
    mem['h65C8]=8'h00; mem['h65C9]=8'h00; mem['h65CA]=8'h00; mem['h65CB]=8'h00;
    mem['h65CC]=8'h00; mem['h65CD]=8'h00; mem['h65CE]=8'h00; mem['h65CF]=8'h00;
    mem['h65D0]=8'h00; mem['h65D1]=8'h00; mem['h65D2]=8'h00; mem['h65D3]=8'h00;
    mem['h65D4]=8'h00; mem['h65D5]=8'h00; mem['h65D6]=8'h00; mem['h65D7]=8'h00;
    mem['h65D8]=8'h00; mem['h65D9]=8'h00; mem['h65DA]=8'h00; mem['h65DB]=8'h00;
    mem['h65DC]=8'h00; mem['h65DD]=8'h00; mem['h65DE]=8'h00; mem['h65DF]=8'h00;
    mem['h65E0]=8'h00; mem['h65E1]=8'h00; mem['h65E2]=8'h00; mem['h65E3]=8'h00;
    mem['h65E4]=8'h00; mem['h65E5]=8'h00; mem['h65E6]=8'h00; mem['h65E7]=8'h00;
    mem['h65E8]=8'h00; mem['h65E9]=8'h00; mem['h65EA]=8'h00; mem['h65EB]=8'h00;
    mem['h65EC]=8'h00; mem['h65ED]=8'h00; mem['h65EE]=8'h00; mem['h65EF]=8'h00;
    mem['h65F0]=8'h00; mem['h65F1]=8'h00; mem['h65F2]=8'h00; mem['h65F3]=8'h00;
    mem['h65F4]=8'h00; mem['h65F5]=8'h00; mem['h65F6]=8'h00; mem['h65F7]=8'h00;
    mem['h65F8]=8'h00; mem['h65F9]=8'h00; mem['h65FA]=8'h00; mem['h65FB]=8'h00;
    mem['h65FC]=8'h00; mem['h65FD]=8'h00; mem['h65FE]=8'h00; mem['h65FF]=8'h00;
    mem['h6600]=8'h00; mem['h6601]=8'h00; mem['h6602]=8'h00; mem['h6603]=8'h00;
    mem['h6604]=8'h00; mem['h6605]=8'h00; mem['h6606]=8'h00; mem['h6607]=8'h00;
    mem['h6608]=8'h00; mem['h6609]=8'h00; mem['h660A]=8'h00; mem['h660B]=8'h00;
    mem['h660C]=8'h00; mem['h660D]=8'h00; mem['h660E]=8'h00; mem['h660F]=8'h00;
    mem['h6610]=8'h00; mem['h6611]=8'h00; mem['h6612]=8'h00; mem['h6613]=8'h00;
    mem['h6614]=8'h00; mem['h6615]=8'h00; mem['h6616]=8'h00; mem['h6617]=8'h00;
    mem['h6618]=8'h00; mem['h6619]=8'h00; mem['h661A]=8'h00; mem['h661B]=8'h00;
    mem['h661C]=8'h00; mem['h661D]=8'h00; mem['h661E]=8'h00; mem['h661F]=8'h00;
    mem['h6620]=8'h00; mem['h6621]=8'h00; mem['h6622]=8'h00; mem['h6623]=8'h00;
    mem['h6624]=8'h00; mem['h6625]=8'h00; mem['h6626]=8'h00; mem['h6627]=8'h00;
    mem['h6628]=8'h00; mem['h6629]=8'h00; mem['h662A]=8'h00; mem['h662B]=8'h00;
    mem['h662C]=8'h00; mem['h662D]=8'h00; mem['h662E]=8'h00; mem['h662F]=8'h00;
    mem['h6630]=8'h00; mem['h6631]=8'h00; mem['h6632]=8'h00; mem['h6633]=8'h00;
    mem['h6634]=8'h00; mem['h6635]=8'h00; mem['h6636]=8'h00; mem['h6637]=8'h00;
    mem['h6638]=8'h00; mem['h6639]=8'h00; mem['h663A]=8'h00; mem['h663B]=8'h00;
    mem['h663C]=8'h00; mem['h663D]=8'h00; mem['h663E]=8'h00; mem['h663F]=8'h00;
    mem['h6640]=8'h00; mem['h6641]=8'h00; mem['h6642]=8'h00; mem['h6643]=8'h00;
    mem['h6644]=8'h00; mem['h6645]=8'h00; mem['h6646]=8'h00; mem['h6647]=8'h00;
    mem['h6648]=8'h00; mem['h6649]=8'h00; mem['h664A]=8'h00; mem['h664B]=8'h00;
    mem['h664C]=8'h00; mem['h664D]=8'h00; mem['h664E]=8'h00; mem['h664F]=8'h00;
    mem['h6650]=8'h00; mem['h6651]=8'h00; mem['h6652]=8'h00; mem['h6653]=8'h00;
    mem['h6654]=8'h00; mem['h6655]=8'h00; mem['h6656]=8'h00; mem['h6657]=8'h00;
    mem['h6658]=8'h00; mem['h6659]=8'h00; mem['h665A]=8'h00; mem['h665B]=8'h00;
    mem['h665C]=8'h00; mem['h665D]=8'h00; mem['h665E]=8'h00; mem['h665F]=8'h00;
    mem['h6660]=8'h00; mem['h6661]=8'h00; mem['h6662]=8'h00; mem['h6663]=8'h00;
    mem['h6664]=8'h00; mem['h6665]=8'h00; mem['h6666]=8'h00; mem['h6667]=8'h00;
    mem['h6668]=8'h00; mem['h6669]=8'h00; mem['h666A]=8'h00; mem['h666B]=8'h00;
    mem['h666C]=8'h00; mem['h666D]=8'h00; mem['h666E]=8'h00; mem['h666F]=8'h00;
    mem['h6670]=8'h00; mem['h6671]=8'h00; mem['h6672]=8'h00; mem['h6673]=8'h00;
    mem['h6674]=8'h00; mem['h6675]=8'h00; mem['h6676]=8'h00; mem['h6677]=8'h00;
    mem['h6678]=8'h00; mem['h6679]=8'h00; mem['h667A]=8'h00; mem['h667B]=8'h00;
    mem['h667C]=8'h00; mem['h667D]=8'h00; mem['h667E]=8'h00; mem['h667F]=8'h00;
    mem['h6680]=8'h00; mem['h6681]=8'h00; mem['h6682]=8'h00; mem['h6683]=8'h00;
    mem['h6684]=8'h00; mem['h6685]=8'h00; mem['h6686]=8'h00; mem['h6687]=8'h00;
    mem['h6688]=8'h00; mem['h6689]=8'h00; mem['h668A]=8'h00; mem['h668B]=8'h00;
    mem['h668C]=8'h00; mem['h668D]=8'h00; mem['h668E]=8'h00; mem['h668F]=8'h00;
    mem['h6690]=8'h00; mem['h6691]=8'h00; mem['h6692]=8'h00; mem['h6693]=8'h00;
    mem['h6694]=8'h00; mem['h6695]=8'h00; mem['h6696]=8'h00; mem['h6697]=8'h00;
    mem['h6698]=8'h00; mem['h6699]=8'h00; mem['h669A]=8'h00; mem['h669B]=8'h00;
    mem['h669C]=8'h00; mem['h669D]=8'h00; mem['h669E]=8'h00; mem['h669F]=8'h00;
    mem['h66A0]=8'h00; mem['h66A1]=8'h00; mem['h66A2]=8'h00; mem['h66A3]=8'h00;
    mem['h66A4]=8'h00; mem['h66A5]=8'h00; mem['h66A6]=8'h00; mem['h66A7]=8'h00;
    mem['h66A8]=8'h00; mem['h66A9]=8'h00; mem['h66AA]=8'h00; mem['h66AB]=8'h00;
    mem['h66AC]=8'h00; mem['h66AD]=8'h00; mem['h66AE]=8'h00; mem['h66AF]=8'h00;
    mem['h66B0]=8'h00; mem['h66B1]=8'h00; mem['h66B2]=8'h00; mem['h66B3]=8'h00;
    mem['h66B4]=8'h00; mem['h66B5]=8'h00; mem['h66B6]=8'h00; mem['h66B7]=8'h00;
    mem['h66B8]=8'h00; mem['h66B9]=8'h00; mem['h66BA]=8'h00; mem['h66BB]=8'h00;
    mem['h66BC]=8'h00; mem['h66BD]=8'h00; mem['h66BE]=8'h00; mem['h66BF]=8'h00;
    mem['h66C0]=8'h00; mem['h66C1]=8'h00; mem['h66C2]=8'h00; mem['h66C3]=8'h00;
    mem['h66C4]=8'h00; mem['h66C5]=8'h00; mem['h66C6]=8'h00; mem['h66C7]=8'h00;
    mem['h66C8]=8'h00; mem['h66C9]=8'h00; mem['h66CA]=8'h00; mem['h66CB]=8'h00;
    mem['h66CC]=8'h00; mem['h66CD]=8'h00; mem['h66CE]=8'h00; mem['h66CF]=8'h00;
    mem['h66D0]=8'h00; mem['h66D1]=8'h00; mem['h66D2]=8'h00; mem['h66D3]=8'h00;
    mem['h66D4]=8'h00; mem['h66D5]=8'h00; mem['h66D6]=8'h00; mem['h66D7]=8'h00;
    mem['h66D8]=8'h00; mem['h66D9]=8'h00; mem['h66DA]=8'h00; mem['h66DB]=8'h00;
    mem['h66DC]=8'h00; mem['h66DD]=8'h00; mem['h66DE]=8'h00; mem['h66DF]=8'h00;
    mem['h66E0]=8'h00; mem['h66E1]=8'h00; mem['h66E2]=8'h00; mem['h66E3]=8'h00;
    mem['h66E4]=8'h00; mem['h66E5]=8'h00; mem['h66E6]=8'h00; mem['h66E7]=8'h00;
    mem['h66E8]=8'h00; mem['h66E9]=8'h00; mem['h66EA]=8'h00; mem['h66EB]=8'h00;
    mem['h66EC]=8'h00; mem['h66ED]=8'h00; mem['h66EE]=8'h00; mem['h66EF]=8'h00;
    mem['h66F0]=8'h00; mem['h66F1]=8'h00; mem['h66F2]=8'h00; mem['h66F3]=8'h00;
    mem['h66F4]=8'h00; mem['h66F5]=8'h00; mem['h66F6]=8'h00; mem['h66F7]=8'h00;
    mem['h66F8]=8'h00; mem['h66F9]=8'h00; mem['h66FA]=8'h00; mem['h66FB]=8'h00;
    mem['h66FC]=8'h00; mem['h66FD]=8'h00; mem['h66FE]=8'h00; mem['h66FF]=8'h00;
    mem['h6700]=8'h00; mem['h6701]=8'h00; mem['h6702]=8'h00; mem['h6703]=8'h00;
    mem['h6704]=8'h00; mem['h6705]=8'h00; mem['h6706]=8'h00; mem['h6707]=8'h00;
    mem['h6708]=8'h00; mem['h6709]=8'h00; mem['h670A]=8'h00; mem['h670B]=8'h00;
    mem['h670C]=8'h00; mem['h670D]=8'h00; mem['h670E]=8'h00; mem['h670F]=8'h00;
    mem['h6710]=8'h00; mem['h6711]=8'h00; mem['h6712]=8'h00; mem['h6713]=8'h00;
    mem['h6714]=8'h00; mem['h6715]=8'h00; mem['h6716]=8'h00; mem['h6717]=8'h00;
    mem['h6718]=8'h00; mem['h6719]=8'h00; mem['h671A]=8'h00; mem['h671B]=8'h00;
    mem['h671C]=8'h00; mem['h671D]=8'h00; mem['h671E]=8'h00; mem['h671F]=8'h00;
    mem['h6720]=8'h00; mem['h6721]=8'h00; mem['h6722]=8'h00; mem['h6723]=8'h00;
    mem['h6724]=8'h00; mem['h6725]=8'h00; mem['h6726]=8'h00; mem['h6727]=8'h00;
    mem['h6728]=8'h00; mem['h6729]=8'h00; mem['h672A]=8'h00; mem['h672B]=8'h00;
    mem['h672C]=8'h00; mem['h672D]=8'h00; mem['h672E]=8'h00; mem['h672F]=8'h00;
    mem['h6730]=8'h00; mem['h6731]=8'h00; mem['h6732]=8'h00; mem['h6733]=8'h00;
    mem['h6734]=8'h00; mem['h6735]=8'h00; mem['h6736]=8'h00; mem['h6737]=8'h00;
    mem['h6738]=8'h00; mem['h6739]=8'h00; mem['h673A]=8'h00; mem['h673B]=8'h00;
    mem['h673C]=8'h00; mem['h673D]=8'h00; mem['h673E]=8'h00; mem['h673F]=8'h00;
    mem['h6740]=8'h00; mem['h6741]=8'h00; mem['h6742]=8'h00; mem['h6743]=8'h00;
    mem['h6744]=8'h00; mem['h6745]=8'h00; mem['h6746]=8'h00; mem['h6747]=8'h00;
    mem['h6748]=8'h00; mem['h6749]=8'h00; mem['h674A]=8'h00; mem['h674B]=8'h00;
    mem['h674C]=8'h00; mem['h674D]=8'h00; mem['h674E]=8'h00; mem['h674F]=8'h00;
    mem['h6750]=8'h00; mem['h6751]=8'h00; mem['h6752]=8'h00; mem['h6753]=8'h00;
    mem['h6754]=8'h00; mem['h6755]=8'h00; mem['h6756]=8'h00; mem['h6757]=8'h00;
    mem['h6758]=8'h00; mem['h6759]=8'h00; mem['h675A]=8'h00; mem['h675B]=8'h00;
    mem['h675C]=8'h00; mem['h675D]=8'h00; mem['h675E]=8'h00; mem['h675F]=8'h00;
    mem['h6760]=8'h00; mem['h6761]=8'h00; mem['h6762]=8'h00; mem['h6763]=8'h00;
    mem['h6764]=8'h00; mem['h6765]=8'h00; mem['h6766]=8'h00; mem['h6767]=8'h00;
    mem['h6768]=8'h00; mem['h6769]=8'h00; mem['h676A]=8'h00; mem['h676B]=8'h00;
    mem['h676C]=8'h00; mem['h676D]=8'h00; mem['h676E]=8'h00; mem['h676F]=8'h00;
    mem['h6770]=8'h00; mem['h6771]=8'h00; mem['h6772]=8'h00; mem['h6773]=8'h00;
    mem['h6774]=8'h00; mem['h6775]=8'h00; mem['h6776]=8'h00; mem['h6777]=8'h00;
    mem['h6778]=8'h00; mem['h6779]=8'h00; mem['h677A]=8'h00; mem['h677B]=8'h00;
    mem['h677C]=8'h00; mem['h677D]=8'h00; mem['h677E]=8'h00; mem['h677F]=8'h00;
    mem['h6780]=8'h00; mem['h6781]=8'h00; mem['h6782]=8'h00; mem['h6783]=8'h00;
    mem['h6784]=8'h00; mem['h6785]=8'h00; mem['h6786]=8'h00; mem['h6787]=8'h00;
    mem['h6788]=8'h00; mem['h6789]=8'h00; mem['h678A]=8'h00; mem['h678B]=8'h00;
    mem['h678C]=8'h00; mem['h678D]=8'h00; mem['h678E]=8'h00; mem['h678F]=8'h00;
    mem['h6790]=8'h00; mem['h6791]=8'h00; mem['h6792]=8'h00; mem['h6793]=8'h00;
    mem['h6794]=8'h00; mem['h6795]=8'h00; mem['h6796]=8'h00; mem['h6797]=8'h00;
    mem['h6798]=8'h00; mem['h6799]=8'h00; mem['h679A]=8'h00; mem['h679B]=8'h00;
    mem['h679C]=8'h00; mem['h679D]=8'h00; mem['h679E]=8'h00; mem['h679F]=8'h00;
    mem['h67A0]=8'h00; mem['h67A1]=8'h00; mem['h67A2]=8'h00; mem['h67A3]=8'h00;
    mem['h67A4]=8'h00; mem['h67A5]=8'h00; mem['h67A6]=8'h00; mem['h67A7]=8'h00;
    mem['h67A8]=8'h00; mem['h67A9]=8'h00; mem['h67AA]=8'h00; mem['h67AB]=8'h00;
    mem['h67AC]=8'h00; mem['h67AD]=8'h00; mem['h67AE]=8'h00; mem['h67AF]=8'h00;
    mem['h67B0]=8'h00; mem['h67B1]=8'h00; mem['h67B2]=8'h00; mem['h67B3]=8'h00;
    mem['h67B4]=8'h00; mem['h67B5]=8'h00; mem['h67B6]=8'h00; mem['h67B7]=8'h00;
    mem['h67B8]=8'h00; mem['h67B9]=8'h00; mem['h67BA]=8'h00; mem['h67BB]=8'h00;
    mem['h67BC]=8'h00; mem['h67BD]=8'h00; mem['h67BE]=8'h00; mem['h67BF]=8'h00;
    mem['h67C0]=8'h00; mem['h67C1]=8'h00; mem['h67C2]=8'h00; mem['h67C3]=8'h00;
    mem['h67C4]=8'h00; mem['h67C5]=8'h00; mem['h67C6]=8'h00; mem['h67C7]=8'h00;
    mem['h67C8]=8'h00; mem['h67C9]=8'h00; mem['h67CA]=8'h00; mem['h67CB]=8'h00;
    mem['h67CC]=8'h00; mem['h67CD]=8'h00; mem['h67CE]=8'h00; mem['h67CF]=8'h00;
    mem['h67D0]=8'h00; mem['h67D1]=8'h00; mem['h67D2]=8'h00; mem['h67D3]=8'h00;
    mem['h67D4]=8'h00; mem['h67D5]=8'h00; mem['h67D6]=8'h00; mem['h67D7]=8'h00;
    mem['h67D8]=8'h00; mem['h67D9]=8'h00; mem['h67DA]=8'h00; mem['h67DB]=8'h00;
    mem['h67DC]=8'h00; mem['h67DD]=8'h00; mem['h67DE]=8'h00; mem['h67DF]=8'h00;
    mem['h67E0]=8'h00; mem['h67E1]=8'h00; mem['h67E2]=8'h00; mem['h67E3]=8'h00;
    mem['h67E4]=8'h00; mem['h67E5]=8'h00; mem['h67E6]=8'h00; mem['h67E7]=8'h00;
    mem['h67E8]=8'h00; mem['h67E9]=8'h00; mem['h67EA]=8'h00; mem['h67EB]=8'h00;
    mem['h67EC]=8'h00; mem['h67ED]=8'h00; mem['h67EE]=8'h00; mem['h67EF]=8'h00;
    mem['h67F0]=8'h00; mem['h67F1]=8'h00; mem['h67F2]=8'h00; mem['h67F3]=8'h00;
    mem['h67F4]=8'h00; mem['h67F5]=8'h00; mem['h67F6]=8'h00; mem['h67F7]=8'h00;
    mem['h67F8]=8'h00; mem['h67F9]=8'h00; mem['h67FA]=8'h00; mem['h67FB]=8'h00;
    mem['h67FC]=8'h00; mem['h67FD]=8'h00; mem['h67FE]=8'h00; mem['h67FF]=8'h00;
    mem['h6800]=8'h00; mem['h6801]=8'h00; mem['h6802]=8'h00; mem['h6803]=8'h00;
    mem['h6804]=8'h00; mem['h6805]=8'h00; mem['h6806]=8'h00; mem['h6807]=8'h00;
    mem['h6808]=8'h00; mem['h6809]=8'h00; mem['h680A]=8'h00; mem['h680B]=8'h00;
    mem['h680C]=8'h00; mem['h680D]=8'h00; mem['h680E]=8'h00; mem['h680F]=8'h00;
    mem['h6810]=8'h00; mem['h6811]=8'h00; mem['h6812]=8'h00; mem['h6813]=8'h00;
    mem['h6814]=8'h00; mem['h6815]=8'h00; mem['h6816]=8'h00; mem['h6817]=8'h00;
    mem['h6818]=8'h00; mem['h6819]=8'h00; mem['h681A]=8'h00; mem['h681B]=8'h00;
    mem['h681C]=8'h00; mem['h681D]=8'h00; mem['h681E]=8'h00; mem['h681F]=8'h00;
    mem['h6820]=8'h00; mem['h6821]=8'h00; mem['h6822]=8'h00; mem['h6823]=8'h00;
    mem['h6824]=8'h00; mem['h6825]=8'h00; mem['h6826]=8'h00; mem['h6827]=8'h00;
    mem['h6828]=8'h00; mem['h6829]=8'h00; mem['h682A]=8'h00; mem['h682B]=8'h00;
    mem['h682C]=8'h00; mem['h682D]=8'h00; mem['h682E]=8'h00; mem['h682F]=8'h00;
    mem['h6830]=8'h00; mem['h6831]=8'h00; mem['h6832]=8'h00; mem['h6833]=8'h00;
    mem['h6834]=8'h00; mem['h6835]=8'h00; mem['h6836]=8'h00; mem['h6837]=8'h00;
    mem['h6838]=8'h00; mem['h6839]=8'h00; mem['h683A]=8'h00; mem['h683B]=8'h00;
    mem['h683C]=8'h00; mem['h683D]=8'h00; mem['h683E]=8'h00; mem['h683F]=8'h00;
    mem['h6840]=8'h00; mem['h6841]=8'h00; mem['h6842]=8'h00; mem['h6843]=8'h00;
    mem['h6844]=8'h00; mem['h6845]=8'h00; mem['h6846]=8'h00; mem['h6847]=8'h00;
    mem['h6848]=8'h00; mem['h6849]=8'h00; mem['h684A]=8'h00; mem['h684B]=8'h00;
    mem['h684C]=8'h00; mem['h684D]=8'h00; mem['h684E]=8'h00; mem['h684F]=8'h00;
    mem['h6850]=8'h00; mem['h6851]=8'h00; mem['h6852]=8'h00; mem['h6853]=8'h00;
    mem['h6854]=8'h00; mem['h6855]=8'h00; mem['h6856]=8'h00; mem['h6857]=8'h00;
    mem['h6858]=8'h00; mem['h6859]=8'h00; mem['h685A]=8'h00; mem['h685B]=8'h00;
    mem['h685C]=8'h00; mem['h685D]=8'h00; mem['h685E]=8'h00; mem['h685F]=8'h00;
    mem['h6860]=8'h00; mem['h6861]=8'h00; mem['h6862]=8'h00; mem['h6863]=8'h00;
    mem['h6864]=8'h00; mem['h6865]=8'h00; mem['h6866]=8'h00; mem['h6867]=8'h00;
    mem['h6868]=8'h00; mem['h6869]=8'h00; mem['h686A]=8'h00; mem['h686B]=8'h00;
    mem['h686C]=8'h00; mem['h686D]=8'h00; mem['h686E]=8'h00; mem['h686F]=8'h00;
    mem['h6870]=8'h00; mem['h6871]=8'h00; mem['h6872]=8'h00; mem['h6873]=8'h00;
    mem['h6874]=8'h00; mem['h6875]=8'h00; mem['h6876]=8'h00; mem['h6877]=8'h00;
    mem['h6878]=8'h00; mem['h6879]=8'h00; mem['h687A]=8'h00; mem['h687B]=8'h00;
    mem['h687C]=8'h00; mem['h687D]=8'h00; mem['h687E]=8'h00; mem['h687F]=8'h00;
    mem['h6880]=8'h00; mem['h6881]=8'h00; mem['h6882]=8'h00; mem['h6883]=8'h00;
    mem['h6884]=8'h00; mem['h6885]=8'h00; mem['h6886]=8'h00; mem['h6887]=8'h00;
    mem['h6888]=8'h00; mem['h6889]=8'h00; mem['h688A]=8'h00; mem['h688B]=8'h00;
    mem['h688C]=8'h00; mem['h688D]=8'h00; mem['h688E]=8'h00; mem['h688F]=8'h00;
    mem['h6890]=8'h00; mem['h6891]=8'h00; mem['h6892]=8'h00; mem['h6893]=8'h00;
    mem['h6894]=8'h00; mem['h6895]=8'h00; mem['h6896]=8'h00; mem['h6897]=8'h00;
    mem['h6898]=8'h00; mem['h6899]=8'h00; mem['h689A]=8'h00; mem['h689B]=8'h00;
    mem['h689C]=8'h00; mem['h689D]=8'h00; mem['h689E]=8'h00; mem['h689F]=8'h00;
    mem['h68A0]=8'h00; mem['h68A1]=8'h00; mem['h68A2]=8'h00; mem['h68A3]=8'h00;
    mem['h68A4]=8'h00; mem['h68A5]=8'h00; mem['h68A6]=8'h00; mem['h68A7]=8'h00;
    mem['h68A8]=8'h00; mem['h68A9]=8'h00; mem['h68AA]=8'h00; mem['h68AB]=8'h00;
    mem['h68AC]=8'h00; mem['h68AD]=8'h00; mem['h68AE]=8'h00; mem['h68AF]=8'h00;
    mem['h68B0]=8'h00; mem['h68B1]=8'h00; mem['h68B2]=8'h00; mem['h68B3]=8'h00;
    mem['h68B4]=8'h00; mem['h68B5]=8'h00; mem['h68B6]=8'h00; mem['h68B7]=8'h00;
    mem['h68B8]=8'h00; mem['h68B9]=8'h00; mem['h68BA]=8'h00; mem['h68BB]=8'h00;
    mem['h68BC]=8'h00; mem['h68BD]=8'h00; mem['h68BE]=8'h00; mem['h68BF]=8'h00;
    mem['h68C0]=8'h00; mem['h68C1]=8'h00; mem['h68C2]=8'h00; mem['h68C3]=8'h00;
    mem['h68C4]=8'h00; mem['h68C5]=8'h00; mem['h68C6]=8'h00; mem['h68C7]=8'h00;
    mem['h68C8]=8'h00; mem['h68C9]=8'h00; mem['h68CA]=8'h00; mem['h68CB]=8'h00;
    mem['h68CC]=8'h00; mem['h68CD]=8'h00; mem['h68CE]=8'h00; mem['h68CF]=8'h00;
    mem['h68D0]=8'h00; mem['h68D1]=8'h00; mem['h68D2]=8'h00; mem['h68D3]=8'h00;
    mem['h68D4]=8'h00; mem['h68D5]=8'h00; mem['h68D6]=8'h00; mem['h68D7]=8'h00;
    mem['h68D8]=8'h00; mem['h68D9]=8'h00; mem['h68DA]=8'h00; mem['h68DB]=8'h00;
    mem['h68DC]=8'h00; mem['h68DD]=8'h00; mem['h68DE]=8'h00; mem['h68DF]=8'h00;
    mem['h68E0]=8'h00; mem['h68E1]=8'h00; mem['h68E2]=8'h00; mem['h68E3]=8'h00;
    mem['h68E4]=8'h00; mem['h68E5]=8'h00; mem['h68E6]=8'h00; mem['h68E7]=8'h00;
    mem['h68E8]=8'h00; mem['h68E9]=8'h00; mem['h68EA]=8'h00; mem['h68EB]=8'h00;
    mem['h68EC]=8'h00; mem['h68ED]=8'h00; mem['h68EE]=8'h00; mem['h68EF]=8'h00;
    mem['h68F0]=8'h00; mem['h68F1]=8'h00; mem['h68F2]=8'h00; mem['h68F3]=8'h00;
    mem['h68F4]=8'h00; mem['h68F5]=8'h00; mem['h68F6]=8'h00; mem['h68F7]=8'h00;
    mem['h68F8]=8'h00; mem['h68F9]=8'h00; mem['h68FA]=8'h00; mem['h68FB]=8'h00;
    mem['h68FC]=8'h00; mem['h68FD]=8'h00; mem['h68FE]=8'h00; mem['h68FF]=8'h00;
    mem['h6900]=8'h00; mem['h6901]=8'h00; mem['h6902]=8'h00; mem['h6903]=8'h00;
    mem['h6904]=8'h00; mem['h6905]=8'h00; mem['h6906]=8'h00; mem['h6907]=8'h00;
    mem['h6908]=8'h00; mem['h6909]=8'h00; mem['h690A]=8'h00; mem['h690B]=8'h00;
    mem['h690C]=8'h00; mem['h690D]=8'h00; mem['h690E]=8'h00; mem['h690F]=8'h00;
    mem['h6910]=8'h00; mem['h6911]=8'h00; mem['h6912]=8'h00; mem['h6913]=8'h00;
    mem['h6914]=8'h00; mem['h6915]=8'h00; mem['h6916]=8'h00; mem['h6917]=8'h00;
    mem['h6918]=8'h00; mem['h6919]=8'h00; mem['h691A]=8'h00; mem['h691B]=8'h00;
    mem['h691C]=8'h00; mem['h691D]=8'h00; mem['h691E]=8'h00; mem['h691F]=8'h00;
    mem['h6920]=8'h00; mem['h6921]=8'h00; mem['h6922]=8'h00; mem['h6923]=8'h00;
    mem['h6924]=8'h00; mem['h6925]=8'h00; mem['h6926]=8'h00; mem['h6927]=8'h00;
    mem['h6928]=8'h00; mem['h6929]=8'h00; mem['h692A]=8'h00; mem['h692B]=8'h00;
    mem['h692C]=8'h00; mem['h692D]=8'h00; mem['h692E]=8'h00; mem['h692F]=8'h00;
    mem['h6930]=8'h00; mem['h6931]=8'h00; mem['h6932]=8'h00; mem['h6933]=8'h00;
    mem['h6934]=8'h00; mem['h6935]=8'h00; mem['h6936]=8'h00; mem['h6937]=8'h00;
    mem['h6938]=8'h00; mem['h6939]=8'h00; mem['h693A]=8'h00; mem['h693B]=8'h00;
    mem['h693C]=8'h00; mem['h693D]=8'h00; mem['h693E]=8'h00; mem['h693F]=8'h00;
    mem['h6940]=8'h00; mem['h6941]=8'h00; mem['h6942]=8'h00; mem['h6943]=8'h00;
    mem['h6944]=8'h00; mem['h6945]=8'h00; mem['h6946]=8'h00; mem['h6947]=8'h00;
    mem['h6948]=8'h00; mem['h6949]=8'h00; mem['h694A]=8'h00; mem['h694B]=8'h00;
    mem['h694C]=8'h00; mem['h694D]=8'h00; mem['h694E]=8'h00; mem['h694F]=8'h00;
    mem['h6950]=8'h00; mem['h6951]=8'h00; mem['h6952]=8'h00; mem['h6953]=8'h00;
    mem['h6954]=8'h00; mem['h6955]=8'h00; mem['h6956]=8'h00; mem['h6957]=8'h00;
    mem['h6958]=8'h00; mem['h6959]=8'h00; mem['h695A]=8'h00; mem['h695B]=8'h00;
    mem['h695C]=8'h00; mem['h695D]=8'h00; mem['h695E]=8'h00; mem['h695F]=8'h00;
    mem['h6960]=8'h00; mem['h6961]=8'h00; mem['h6962]=8'h00; mem['h6963]=8'h00;
    mem['h6964]=8'h00; mem['h6965]=8'h00; mem['h6966]=8'h00; mem['h6967]=8'h00;
    mem['h6968]=8'h00; mem['h6969]=8'h00; mem['h696A]=8'h00; mem['h696B]=8'h00;
    mem['h696C]=8'h00; mem['h696D]=8'h00; mem['h696E]=8'h00; mem['h696F]=8'h00;
    mem['h6970]=8'h00; mem['h6971]=8'h00; mem['h6972]=8'h00; mem['h6973]=8'h00;
    mem['h6974]=8'h00; mem['h6975]=8'h00; mem['h6976]=8'h00; mem['h6977]=8'h00;
    mem['h6978]=8'h00; mem['h6979]=8'h00; mem['h697A]=8'h00; mem['h697B]=8'h00;
    mem['h697C]=8'h00; mem['h697D]=8'h00; mem['h697E]=8'h00; mem['h697F]=8'h00;
    mem['h6980]=8'h00; mem['h6981]=8'h00; mem['h6982]=8'h00; mem['h6983]=8'h00;
    mem['h6984]=8'h00; mem['h6985]=8'h00; mem['h6986]=8'h00; mem['h6987]=8'h00;
    mem['h6988]=8'h00; mem['h6989]=8'h00; mem['h698A]=8'h00; mem['h698B]=8'h00;
    mem['h698C]=8'h00; mem['h698D]=8'h00; mem['h698E]=8'h00; mem['h698F]=8'h00;
    mem['h6990]=8'h00; mem['h6991]=8'h00; mem['h6992]=8'h00; mem['h6993]=8'h00;
    mem['h6994]=8'h00; mem['h6995]=8'h00; mem['h6996]=8'h00; mem['h6997]=8'h00;
    mem['h6998]=8'h00; mem['h6999]=8'h00; mem['h699A]=8'h00; mem['h699B]=8'h00;
    mem['h699C]=8'h00; mem['h699D]=8'h00; mem['h699E]=8'h00; mem['h699F]=8'h00;
    mem['h69A0]=8'h00; mem['h69A1]=8'h00; mem['h69A2]=8'h00; mem['h69A3]=8'h00;
    mem['h69A4]=8'h00; mem['h69A5]=8'h00; mem['h69A6]=8'h00; mem['h69A7]=8'h00;
    mem['h69A8]=8'h00; mem['h69A9]=8'h00; mem['h69AA]=8'h00; mem['h69AB]=8'h00;
    mem['h69AC]=8'h00; mem['h69AD]=8'h00; mem['h69AE]=8'h00; mem['h69AF]=8'h00;
    mem['h69B0]=8'h00; mem['h69B1]=8'h00; mem['h69B2]=8'h00; mem['h69B3]=8'h00;
    mem['h69B4]=8'h00; mem['h69B5]=8'h00; mem['h69B6]=8'h00; mem['h69B7]=8'h00;
    mem['h69B8]=8'h00; mem['h69B9]=8'h00; mem['h69BA]=8'h00; mem['h69BB]=8'h00;
    mem['h69BC]=8'h00; mem['h69BD]=8'h00; mem['h69BE]=8'h00; mem['h69BF]=8'h00;
    mem['h69C0]=8'h00; mem['h69C1]=8'h00; mem['h69C2]=8'h00; mem['h69C3]=8'h00;
    mem['h69C4]=8'h00; mem['h69C5]=8'h00; mem['h69C6]=8'h00; mem['h69C7]=8'h00;
    mem['h69C8]=8'h00; mem['h69C9]=8'h00; mem['h69CA]=8'h00; mem['h69CB]=8'h00;
    mem['h69CC]=8'h00; mem['h69CD]=8'h00; mem['h69CE]=8'h00; mem['h69CF]=8'h00;
    mem['h69D0]=8'h00; mem['h69D1]=8'h00; mem['h69D2]=8'h00; mem['h69D3]=8'h00;
    mem['h69D4]=8'h00; mem['h69D5]=8'h00; mem['h69D6]=8'h00; mem['h69D7]=8'h00;
    mem['h69D8]=8'h00; mem['h69D9]=8'h00; mem['h69DA]=8'h00; mem['h69DB]=8'h00;
    mem['h69DC]=8'h00; mem['h69DD]=8'h00; mem['h69DE]=8'h00; mem['h69DF]=8'h00;
    mem['h69E0]=8'h00; mem['h69E1]=8'h00; mem['h69E2]=8'h00; mem['h69E3]=8'h00;
    mem['h69E4]=8'h00; mem['h69E5]=8'h00; mem['h69E6]=8'h00; mem['h69E7]=8'h00;
    mem['h69E8]=8'h00; mem['h69E9]=8'h00; mem['h69EA]=8'h00; mem['h69EB]=8'h00;
    mem['h69EC]=8'h00; mem['h69ED]=8'h00; mem['h69EE]=8'h00; mem['h69EF]=8'h00;
    mem['h69F0]=8'h00; mem['h69F1]=8'h00; mem['h69F2]=8'h00; mem['h69F3]=8'h00;
    mem['h69F4]=8'h00; mem['h69F5]=8'h00; mem['h69F6]=8'h00; mem['h69F7]=8'h00;
    mem['h69F8]=8'h00; mem['h69F9]=8'h00; mem['h69FA]=8'h00; mem['h69FB]=8'h00;
    mem['h69FC]=8'h00; mem['h69FD]=8'h00; mem['h69FE]=8'h00; mem['h69FF]=8'h00;
    mem['h6A00]=8'h00; mem['h6A01]=8'h00; mem['h6A02]=8'h00; mem['h6A03]=8'h00;
    mem['h6A04]=8'h00; mem['h6A05]=8'h00; mem['h6A06]=8'h00; mem['h6A07]=8'h00;
    mem['h6A08]=8'h00; mem['h6A09]=8'h00; mem['h6A0A]=8'h00; mem['h6A0B]=8'h00;
    mem['h6A0C]=8'h00; mem['h6A0D]=8'h00; mem['h6A0E]=8'h00; mem['h6A0F]=8'h00;
    mem['h6A10]=8'h00; mem['h6A11]=8'h00; mem['h6A12]=8'h00; mem['h6A13]=8'h00;
    mem['h6A14]=8'h00; mem['h6A15]=8'h00; mem['h6A16]=8'h00; mem['h6A17]=8'h00;
    mem['h6A18]=8'h00; mem['h6A19]=8'h00; mem['h6A1A]=8'h00; mem['h6A1B]=8'h00;
    mem['h6A1C]=8'h00; mem['h6A1D]=8'h00; mem['h6A1E]=8'h00; mem['h6A1F]=8'h00;
    mem['h6A20]=8'h00; mem['h6A21]=8'h00; mem['h6A22]=8'h00; mem['h6A23]=8'h00;
    mem['h6A24]=8'h00; mem['h6A25]=8'h00; mem['h6A26]=8'h00; mem['h6A27]=8'h00;
    mem['h6A28]=8'h00; mem['h6A29]=8'h00; mem['h6A2A]=8'h00; mem['h6A2B]=8'h00;
    mem['h6A2C]=8'h00; mem['h6A2D]=8'h00; mem['h6A2E]=8'h00; mem['h6A2F]=8'h00;
    mem['h6A30]=8'h00; mem['h6A31]=8'h00; mem['h6A32]=8'h00; mem['h6A33]=8'h00;
    mem['h6A34]=8'h00; mem['h6A35]=8'h00; mem['h6A36]=8'h00; mem['h6A37]=8'h00;
    mem['h6A38]=8'h00; mem['h6A39]=8'h00; mem['h6A3A]=8'h00; mem['h6A3B]=8'h00;
    mem['h6A3C]=8'h00; mem['h6A3D]=8'h00; mem['h6A3E]=8'h00; mem['h6A3F]=8'h00;
    mem['h6A40]=8'h00; mem['h6A41]=8'h00; mem['h6A42]=8'h00; mem['h6A43]=8'h00;
    mem['h6A44]=8'h00; mem['h6A45]=8'h00; mem['h6A46]=8'h00; mem['h6A47]=8'h00;
    mem['h6A48]=8'h00; mem['h6A49]=8'h00; mem['h6A4A]=8'h00; mem['h6A4B]=8'h00;
    mem['h6A4C]=8'h00; mem['h6A4D]=8'h00; mem['h6A4E]=8'h00; mem['h6A4F]=8'h00;
    mem['h6A50]=8'h00; mem['h6A51]=8'h00; mem['h6A52]=8'h00; mem['h6A53]=8'h00;
    mem['h6A54]=8'h00; mem['h6A55]=8'h00; mem['h6A56]=8'h00; mem['h6A57]=8'h00;
    mem['h6A58]=8'h00; mem['h6A59]=8'h00; mem['h6A5A]=8'h00; mem['h6A5B]=8'h00;
    mem['h6A5C]=8'h00; mem['h6A5D]=8'h00; mem['h6A5E]=8'h00; mem['h6A5F]=8'h00;
    mem['h6A60]=8'h00; mem['h6A61]=8'h00; mem['h6A62]=8'h00; mem['h6A63]=8'h00;
    mem['h6A64]=8'h00; mem['h6A65]=8'h00; mem['h6A66]=8'h00; mem['h6A67]=8'h00;
    mem['h6A68]=8'h00; mem['h6A69]=8'h00; mem['h6A6A]=8'h00; mem['h6A6B]=8'h00;
    mem['h6A6C]=8'h00; mem['h6A6D]=8'h00; mem['h6A6E]=8'h00; mem['h6A6F]=8'h00;
    mem['h6A70]=8'h00; mem['h6A71]=8'h00; mem['h6A72]=8'h00; mem['h6A73]=8'h00;
    mem['h6A74]=8'h00; mem['h6A75]=8'h00; mem['h6A76]=8'h00; mem['h6A77]=8'h00;
    mem['h6A78]=8'h00; mem['h6A79]=8'h00; mem['h6A7A]=8'h00; mem['h6A7B]=8'h00;
    mem['h6A7C]=8'h00; mem['h6A7D]=8'h00; mem['h6A7E]=8'h00; mem['h6A7F]=8'h00;
    mem['h6A80]=8'h00; mem['h6A81]=8'h00; mem['h6A82]=8'h00; mem['h6A83]=8'h00;
    mem['h6A84]=8'h00; mem['h6A85]=8'h00; mem['h6A86]=8'h00; mem['h6A87]=8'h00;
    mem['h6A88]=8'h00; mem['h6A89]=8'h00; mem['h6A8A]=8'h00; mem['h6A8B]=8'h00;
    mem['h6A8C]=8'h00; mem['h6A8D]=8'h00; mem['h6A8E]=8'h00; mem['h6A8F]=8'h00;
    mem['h6A90]=8'h00; mem['h6A91]=8'h00; mem['h6A92]=8'h00; mem['h6A93]=8'h00;
    mem['h6A94]=8'h00; mem['h6A95]=8'h00; mem['h6A96]=8'h00; mem['h6A97]=8'h00;
    mem['h6A98]=8'h00; mem['h6A99]=8'h00; mem['h6A9A]=8'h00; mem['h6A9B]=8'h00;
    mem['h6A9C]=8'h00; mem['h6A9D]=8'h00; mem['h6A9E]=8'h00; mem['h6A9F]=8'h00;
    mem['h6AA0]=8'h00; mem['h6AA1]=8'h00; mem['h6AA2]=8'h00; mem['h6AA3]=8'h00;
    mem['h6AA4]=8'h00; mem['h6AA5]=8'h00; mem['h6AA6]=8'h00; mem['h6AA7]=8'h00;
    mem['h6AA8]=8'h00; mem['h6AA9]=8'h00; mem['h6AAA]=8'h00; mem['h6AAB]=8'h00;
    mem['h6AAC]=8'h00; mem['h6AAD]=8'h00; mem['h6AAE]=8'h00; mem['h6AAF]=8'h00;
    mem['h6AB0]=8'h00; mem['h6AB1]=8'h00; mem['h6AB2]=8'h00; mem['h6AB3]=8'h00;
    mem['h6AB4]=8'h00; mem['h6AB5]=8'h00; mem['h6AB6]=8'h00; mem['h6AB7]=8'h00;
    mem['h6AB8]=8'h00; mem['h6AB9]=8'h00; mem['h6ABA]=8'h00; mem['h6ABB]=8'h00;
    mem['h6ABC]=8'h00; mem['h6ABD]=8'h00; mem['h6ABE]=8'h00; mem['h6ABF]=8'h00;
    mem['h6AC0]=8'h00; mem['h6AC1]=8'h00; mem['h6AC2]=8'h00; mem['h6AC3]=8'h00;
    mem['h6AC4]=8'h00; mem['h6AC5]=8'h00; mem['h6AC6]=8'h00; mem['h6AC7]=8'h00;
    mem['h6AC8]=8'h00; mem['h6AC9]=8'h00; mem['h6ACA]=8'h00; mem['h6ACB]=8'h00;
    mem['h6ACC]=8'h00; mem['h6ACD]=8'h00; mem['h6ACE]=8'h00; mem['h6ACF]=8'h00;
    mem['h6AD0]=8'h00; mem['h6AD1]=8'h00; mem['h6AD2]=8'h00; mem['h6AD3]=8'h00;
    mem['h6AD4]=8'h00; mem['h6AD5]=8'h00; mem['h6AD6]=8'h00; mem['h6AD7]=8'h00;
    mem['h6AD8]=8'h00; mem['h6AD9]=8'h00; mem['h6ADA]=8'h00; mem['h6ADB]=8'h00;
    mem['h6ADC]=8'h00; mem['h6ADD]=8'h00; mem['h6ADE]=8'h00; mem['h6ADF]=8'h00;
    mem['h6AE0]=8'h00; mem['h6AE1]=8'h00; mem['h6AE2]=8'h00; mem['h6AE3]=8'h00;
    mem['h6AE4]=8'h00; mem['h6AE5]=8'h00; mem['h6AE6]=8'h00; mem['h6AE7]=8'h00;
    mem['h6AE8]=8'h00; mem['h6AE9]=8'h00; mem['h6AEA]=8'h00; mem['h6AEB]=8'h00;
    mem['h6AEC]=8'h00; mem['h6AED]=8'h00; mem['h6AEE]=8'h00; mem['h6AEF]=8'h00;
    mem['h6AF0]=8'h00; mem['h6AF1]=8'h00; mem['h6AF2]=8'h00; mem['h6AF3]=8'h00;
    mem['h6AF4]=8'h00; mem['h6AF5]=8'h00; mem['h6AF6]=8'h00; mem['h6AF7]=8'h00;
    mem['h6AF8]=8'h00; mem['h6AF9]=8'h00; mem['h6AFA]=8'h00; mem['h6AFB]=8'h00;
    mem['h6AFC]=8'h00; mem['h6AFD]=8'h00; mem['h6AFE]=8'h00; mem['h6AFF]=8'h00;
    mem['h6B00]=8'h00; mem['h6B01]=8'h00; mem['h6B02]=8'h00; mem['h6B03]=8'h00;
    mem['h6B04]=8'h00; mem['h6B05]=8'h00; mem['h6B06]=8'h00; mem['h6B07]=8'h00;
    mem['h6B08]=8'h00; mem['h6B09]=8'h00; mem['h6B0A]=8'h00; mem['h6B0B]=8'h00;
    mem['h6B0C]=8'h00; mem['h6B0D]=8'h00; mem['h6B0E]=8'h00; mem['h6B0F]=8'h00;
    mem['h6B10]=8'h00; mem['h6B11]=8'h00; mem['h6B12]=8'h00; mem['h6B13]=8'h00;
    mem['h6B14]=8'h00; mem['h6B15]=8'h00; mem['h6B16]=8'h00; mem['h6B17]=8'h00;
    mem['h6B18]=8'h00; mem['h6B19]=8'h00; mem['h6B1A]=8'h00; mem['h6B1B]=8'h00;
    mem['h6B1C]=8'h00; mem['h6B1D]=8'h00; mem['h6B1E]=8'h00; mem['h6B1F]=8'h00;
    mem['h6B20]=8'h00; mem['h6B21]=8'h00; mem['h6B22]=8'h00; mem['h6B23]=8'h00;
    mem['h6B24]=8'h00; mem['h6B25]=8'h00; mem['h6B26]=8'h00; mem['h6B27]=8'h00;
    mem['h6B28]=8'h00; mem['h6B29]=8'h00; mem['h6B2A]=8'h00; mem['h6B2B]=8'h00;
    mem['h6B2C]=8'h00; mem['h6B2D]=8'h00; mem['h6B2E]=8'h00; mem['h6B2F]=8'h00;
    mem['h6B30]=8'h00; mem['h6B31]=8'h00; mem['h6B32]=8'h00; mem['h6B33]=8'h00;
    mem['h6B34]=8'h00; mem['h6B35]=8'h00; mem['h6B36]=8'h00; mem['h6B37]=8'h00;
    mem['h6B38]=8'h00; mem['h6B39]=8'h00; mem['h6B3A]=8'h00; mem['h6B3B]=8'h00;
    mem['h6B3C]=8'h00; mem['h6B3D]=8'h00; mem['h6B3E]=8'h00; mem['h6B3F]=8'h00;
    mem['h6B40]=8'h00; mem['h6B41]=8'h00; mem['h6B42]=8'h00; mem['h6B43]=8'h00;
    mem['h6B44]=8'h00; mem['h6B45]=8'h00; mem['h6B46]=8'h00; mem['h6B47]=8'h00;
    mem['h6B48]=8'h00; mem['h6B49]=8'h00; mem['h6B4A]=8'h00; mem['h6B4B]=8'h00;
    mem['h6B4C]=8'h00; mem['h6B4D]=8'h00; mem['h6B4E]=8'h00; mem['h6B4F]=8'h00;
    mem['h6B50]=8'h00; mem['h6B51]=8'h00; mem['h6B52]=8'h00; mem['h6B53]=8'h00;
    mem['h6B54]=8'h00; mem['h6B55]=8'h00; mem['h6B56]=8'h00; mem['h6B57]=8'h00;
    mem['h6B58]=8'h00; mem['h6B59]=8'h00; mem['h6B5A]=8'h00; mem['h6B5B]=8'h00;
    mem['h6B5C]=8'h00; mem['h6B5D]=8'h00; mem['h6B5E]=8'h00; mem['h6B5F]=8'h00;
    mem['h6B60]=8'h00; mem['h6B61]=8'h00; mem['h6B62]=8'h00; mem['h6B63]=8'h00;
    mem['h6B64]=8'h00; mem['h6B65]=8'h00; mem['h6B66]=8'h00; mem['h6B67]=8'h00;
    mem['h6B68]=8'h00; mem['h6B69]=8'h00; mem['h6B6A]=8'h00; mem['h6B6B]=8'h00;
    mem['h6B6C]=8'h00; mem['h6B6D]=8'h00; mem['h6B6E]=8'h00; mem['h6B6F]=8'h00;
    mem['h6B70]=8'h00; mem['h6B71]=8'h00; mem['h6B72]=8'h00; mem['h6B73]=8'h00;
    mem['h6B74]=8'h00; mem['h6B75]=8'h00; mem['h6B76]=8'h00; mem['h6B77]=8'h00;
    mem['h6B78]=8'h00; mem['h6B79]=8'h00; mem['h6B7A]=8'h00; mem['h6B7B]=8'h00;
    mem['h6B7C]=8'h00; mem['h6B7D]=8'h00; mem['h6B7E]=8'h00; mem['h6B7F]=8'h00;
    mem['h6B80]=8'h00; mem['h6B81]=8'h00; mem['h6B82]=8'h00; mem['h6B83]=8'h00;
    mem['h6B84]=8'h00; mem['h6B85]=8'h00; mem['h6B86]=8'h00; mem['h6B87]=8'h00;
    mem['h6B88]=8'h00; mem['h6B89]=8'h00; mem['h6B8A]=8'h00; mem['h6B8B]=8'h00;
    mem['h6B8C]=8'h00; mem['h6B8D]=8'h00; mem['h6B8E]=8'h00; mem['h6B8F]=8'h00;
    mem['h6B90]=8'h00; mem['h6B91]=8'h00; mem['h6B92]=8'h00; mem['h6B93]=8'h00;
    mem['h6B94]=8'h00; mem['h6B95]=8'h00; mem['h6B96]=8'h00; mem['h6B97]=8'h00;
    mem['h6B98]=8'h00; mem['h6B99]=8'h00; mem['h6B9A]=8'h00; mem['h6B9B]=8'h00;
    mem['h6B9C]=8'h00; mem['h6B9D]=8'h00; mem['h6B9E]=8'h00; mem['h6B9F]=8'h00;
    mem['h6BA0]=8'h00; mem['h6BA1]=8'h00; mem['h6BA2]=8'h00; mem['h6BA3]=8'h00;
    mem['h6BA4]=8'h00; mem['h6BA5]=8'h00; mem['h6BA6]=8'h00; mem['h6BA7]=8'h00;
    mem['h6BA8]=8'h00; mem['h6BA9]=8'h00; mem['h6BAA]=8'h00; mem['h6BAB]=8'h00;
    mem['h6BAC]=8'h00; mem['h6BAD]=8'h00; mem['h6BAE]=8'h00; mem['h6BAF]=8'h00;
    mem['h6BB0]=8'h00; mem['h6BB1]=8'h00; mem['h6BB2]=8'h00; mem['h6BB3]=8'h00;
    mem['h6BB4]=8'h00; mem['h6BB5]=8'h00; mem['h6BB6]=8'h00; mem['h6BB7]=8'h00;
    mem['h6BB8]=8'h00; mem['h6BB9]=8'h00; mem['h6BBA]=8'h00; mem['h6BBB]=8'h00;
    mem['h6BBC]=8'h00; mem['h6BBD]=8'h00; mem['h6BBE]=8'h00; mem['h6BBF]=8'h00;
    mem['h6BC0]=8'h00; mem['h6BC1]=8'h00; mem['h6BC2]=8'h00; mem['h6BC3]=8'h00;
    mem['h6BC4]=8'h00; mem['h6BC5]=8'h00; mem['h6BC6]=8'h00; mem['h6BC7]=8'h00;
    mem['h6BC8]=8'h00; mem['h6BC9]=8'h00; mem['h6BCA]=8'h00; mem['h6BCB]=8'h00;
    mem['h6BCC]=8'h00; mem['h6BCD]=8'h00; mem['h6BCE]=8'h00; mem['h6BCF]=8'h00;
    mem['h6BD0]=8'h00; mem['h6BD1]=8'h00; mem['h6BD2]=8'h00; mem['h6BD3]=8'h00;
    mem['h6BD4]=8'h00; mem['h6BD5]=8'h00; mem['h6BD6]=8'h00; mem['h6BD7]=8'h00;
    mem['h6BD8]=8'h00; mem['h6BD9]=8'h00; mem['h6BDA]=8'h00; mem['h6BDB]=8'h00;
    mem['h6BDC]=8'h00; mem['h6BDD]=8'h00; mem['h6BDE]=8'h00; mem['h6BDF]=8'h00;
    mem['h6BE0]=8'h00; mem['h6BE1]=8'h00; mem['h6BE2]=8'h00; mem['h6BE3]=8'h00;
    mem['h6BE4]=8'h00; mem['h6BE5]=8'h00; mem['h6BE6]=8'h00; mem['h6BE7]=8'h00;
    mem['h6BE8]=8'h00; mem['h6BE9]=8'h00; mem['h6BEA]=8'h00; mem['h6BEB]=8'h00;
    mem['h6BEC]=8'h00; mem['h6BED]=8'h00; mem['h6BEE]=8'h00; mem['h6BEF]=8'h00;
    mem['h6BF0]=8'h00; mem['h6BF1]=8'h00; mem['h6BF2]=8'h00; mem['h6BF3]=8'h00;
    mem['h6BF4]=8'h00; mem['h6BF5]=8'h00; mem['h6BF6]=8'h00; mem['h6BF7]=8'h00;
    mem['h6BF8]=8'h00; mem['h6BF9]=8'h00; mem['h6BFA]=8'h00; mem['h6BFB]=8'h00;
    mem['h6BFC]=8'h00; mem['h6BFD]=8'h00; mem['h6BFE]=8'h00; mem['h6BFF]=8'h00;
    mem['h6C00]=8'h00; mem['h6C01]=8'h00; mem['h6C02]=8'h00; mem['h6C03]=8'h00;
    mem['h6C04]=8'h00; mem['h6C05]=8'h00; mem['h6C06]=8'h00; mem['h6C07]=8'h00;
    mem['h6C08]=8'h00; mem['h6C09]=8'h00; mem['h6C0A]=8'h00; mem['h6C0B]=8'h00;
    mem['h6C0C]=8'h00; mem['h6C0D]=8'h00; mem['h6C0E]=8'h00; mem['h6C0F]=8'h00;
    mem['h6C10]=8'h00; mem['h6C11]=8'h00; mem['h6C12]=8'h00; mem['h6C13]=8'h00;
    mem['h6C14]=8'h00; mem['h6C15]=8'h00; mem['h6C16]=8'h00; mem['h6C17]=8'h00;
    mem['h6C18]=8'h00; mem['h6C19]=8'h00; mem['h6C1A]=8'h00; mem['h6C1B]=8'h00;
    mem['h6C1C]=8'h00; mem['h6C1D]=8'h00; mem['h6C1E]=8'h00; mem['h6C1F]=8'h00;
    mem['h6C20]=8'h00; mem['h6C21]=8'h00; mem['h6C22]=8'h00; mem['h6C23]=8'h00;
    mem['h6C24]=8'h00; mem['h6C25]=8'h00; mem['h6C26]=8'h00; mem['h6C27]=8'h00;
    mem['h6C28]=8'h00; mem['h6C29]=8'h00; mem['h6C2A]=8'h00; mem['h6C2B]=8'h00;
    mem['h6C2C]=8'h00; mem['h6C2D]=8'h00; mem['h6C2E]=8'h00; mem['h6C2F]=8'h00;
    mem['h6C30]=8'h00; mem['h6C31]=8'h00; mem['h6C32]=8'h00; mem['h6C33]=8'h00;
    mem['h6C34]=8'h00; mem['h6C35]=8'h00; mem['h6C36]=8'h00; mem['h6C37]=8'h00;
    mem['h6C38]=8'h00; mem['h6C39]=8'h00; mem['h6C3A]=8'h00; mem['h6C3B]=8'h00;
    mem['h6C3C]=8'h00; mem['h6C3D]=8'h00; mem['h6C3E]=8'h00; mem['h6C3F]=8'h00;
    mem['h6C40]=8'h00; mem['h6C41]=8'h00; mem['h6C42]=8'h00; mem['h6C43]=8'h00;
    mem['h6C44]=8'h00; mem['h6C45]=8'h00; mem['h6C46]=8'h00; mem['h6C47]=8'h00;
    mem['h6C48]=8'h00; mem['h6C49]=8'h00; mem['h6C4A]=8'h00; mem['h6C4B]=8'h00;
    mem['h6C4C]=8'h00; mem['h6C4D]=8'h00; mem['h6C4E]=8'h00; mem['h6C4F]=8'h00;
    mem['h6C50]=8'h00; mem['h6C51]=8'h00; mem['h6C52]=8'h00; mem['h6C53]=8'h00;
    mem['h6C54]=8'h00; mem['h6C55]=8'h00; mem['h6C56]=8'h00; mem['h6C57]=8'h00;
    mem['h6C58]=8'h00; mem['h6C59]=8'h00; mem['h6C5A]=8'h00; mem['h6C5B]=8'h00;
    mem['h6C5C]=8'h00; mem['h6C5D]=8'h00; mem['h6C5E]=8'h00; mem['h6C5F]=8'h00;
    mem['h6C60]=8'h00; mem['h6C61]=8'h00; mem['h6C62]=8'h00; mem['h6C63]=8'h00;
    mem['h6C64]=8'h00; mem['h6C65]=8'h00; mem['h6C66]=8'h00; mem['h6C67]=8'h00;
    mem['h6C68]=8'h00; mem['h6C69]=8'h00; mem['h6C6A]=8'h00; mem['h6C6B]=8'h00;
    mem['h6C6C]=8'h00; mem['h6C6D]=8'h00; mem['h6C6E]=8'h00; mem['h6C6F]=8'h00;
    mem['h6C70]=8'h00; mem['h6C71]=8'h00; mem['h6C72]=8'h00; mem['h6C73]=8'h00;
    mem['h6C74]=8'h00; mem['h6C75]=8'h00; mem['h6C76]=8'h00; mem['h6C77]=8'h00;
    mem['h6C78]=8'h00; mem['h6C79]=8'h00; mem['h6C7A]=8'h00; mem['h6C7B]=8'h00;
    mem['h6C7C]=8'h00; mem['h6C7D]=8'h00; mem['h6C7E]=8'h00; mem['h6C7F]=8'h00;
    mem['h6C80]=8'h00; mem['h6C81]=8'h00; mem['h6C82]=8'h00; mem['h6C83]=8'h00;
    mem['h6C84]=8'h00; mem['h6C85]=8'h00; mem['h6C86]=8'h00; mem['h6C87]=8'h00;
    mem['h6C88]=8'h00; mem['h6C89]=8'h00; mem['h6C8A]=8'h00; mem['h6C8B]=8'h00;
    mem['h6C8C]=8'h00; mem['h6C8D]=8'h00; mem['h6C8E]=8'h00; mem['h6C8F]=8'h00;
    mem['h6C90]=8'h00; mem['h6C91]=8'h00; mem['h6C92]=8'h00; mem['h6C93]=8'h00;
    mem['h6C94]=8'h00; mem['h6C95]=8'h00; mem['h6C96]=8'h00; mem['h6C97]=8'h00;
    mem['h6C98]=8'h00; mem['h6C99]=8'h00; mem['h6C9A]=8'h00; mem['h6C9B]=8'h00;
    mem['h6C9C]=8'h00; mem['h6C9D]=8'h00; mem['h6C9E]=8'h00; mem['h6C9F]=8'h00;
    mem['h6CA0]=8'h00; mem['h6CA1]=8'h00; mem['h6CA2]=8'h00; mem['h6CA3]=8'h00;
    mem['h6CA4]=8'h00; mem['h6CA5]=8'h00; mem['h6CA6]=8'h00; mem['h6CA7]=8'h00;
    mem['h6CA8]=8'h00; mem['h6CA9]=8'h00; mem['h6CAA]=8'h00; mem['h6CAB]=8'h00;
    mem['h6CAC]=8'h00; mem['h6CAD]=8'h00; mem['h6CAE]=8'h00; mem['h6CAF]=8'h00;
    mem['h6CB0]=8'h00; mem['h6CB1]=8'h00; mem['h6CB2]=8'h00; mem['h6CB3]=8'h00;
    mem['h6CB4]=8'h00; mem['h6CB5]=8'h00; mem['h6CB6]=8'h00; mem['h6CB7]=8'h00;
    mem['h6CB8]=8'h00; mem['h6CB9]=8'h00; mem['h6CBA]=8'h00; mem['h6CBB]=8'h00;
    mem['h6CBC]=8'h00; mem['h6CBD]=8'h00; mem['h6CBE]=8'h00; mem['h6CBF]=8'h00;
    mem['h6CC0]=8'h00; mem['h6CC1]=8'h00; mem['h6CC2]=8'h00; mem['h6CC3]=8'h00;
    mem['h6CC4]=8'h00; mem['h6CC5]=8'h00; mem['h6CC6]=8'h00; mem['h6CC7]=8'h00;
    mem['h6CC8]=8'h00; mem['h6CC9]=8'h00; mem['h6CCA]=8'h00; mem['h6CCB]=8'h00;
    mem['h6CCC]=8'h00; mem['h6CCD]=8'h00; mem['h6CCE]=8'h00; mem['h6CCF]=8'h00;
    mem['h6CD0]=8'h00; mem['h6CD1]=8'h00; mem['h6CD2]=8'h00; mem['h6CD3]=8'h00;
    mem['h6CD4]=8'h00; mem['h6CD5]=8'h00; mem['h6CD6]=8'h00; mem['h6CD7]=8'h00;
    mem['h6CD8]=8'h00; mem['h6CD9]=8'h00; mem['h6CDA]=8'h00; mem['h6CDB]=8'h00;
    mem['h6CDC]=8'h00; mem['h6CDD]=8'h00; mem['h6CDE]=8'h00; mem['h6CDF]=8'h00;
    mem['h6CE0]=8'h00; mem['h6CE1]=8'h00; mem['h6CE2]=8'h00; mem['h6CE3]=8'h00;
    mem['h6CE4]=8'h00; mem['h6CE5]=8'h00; mem['h6CE6]=8'h00; mem['h6CE7]=8'h00;
    mem['h6CE8]=8'h00; mem['h6CE9]=8'h00; mem['h6CEA]=8'h00; mem['h6CEB]=8'h00;
    mem['h6CEC]=8'h00; mem['h6CED]=8'h00; mem['h6CEE]=8'h00; mem['h6CEF]=8'h00;
    mem['h6CF0]=8'h00; mem['h6CF1]=8'h00; mem['h6CF2]=8'h00; mem['h6CF3]=8'h00;
    mem['h6CF4]=8'h00; mem['h6CF5]=8'h00; mem['h6CF6]=8'h00; mem['h6CF7]=8'h00;
    mem['h6CF8]=8'h00; mem['h6CF9]=8'h00; mem['h6CFA]=8'h00; mem['h6CFB]=8'h00;
    mem['h6CFC]=8'h00; mem['h6CFD]=8'h00; mem['h6CFE]=8'h00; mem['h6CFF]=8'h00;
    mem['h6D00]=8'h00; mem['h6D01]=8'h00; mem['h6D02]=8'h00; mem['h6D03]=8'h00;
    mem['h6D04]=8'h00; mem['h6D05]=8'h00; mem['h6D06]=8'h00; mem['h6D07]=8'h00;
    mem['h6D08]=8'h00; mem['h6D09]=8'h00; mem['h6D0A]=8'h00; mem['h6D0B]=8'h00;
    mem['h6D0C]=8'h00; mem['h6D0D]=8'h00; mem['h6D0E]=8'h00; mem['h6D0F]=8'h00;
    mem['h6D10]=8'h00; mem['h6D11]=8'h00; mem['h6D12]=8'h00; mem['h6D13]=8'h00;
    mem['h6D14]=8'h00; mem['h6D15]=8'h00; mem['h6D16]=8'h00; mem['h6D17]=8'h00;
    mem['h6D18]=8'h00; mem['h6D19]=8'h00; mem['h6D1A]=8'h00; mem['h6D1B]=8'h00;
    mem['h6D1C]=8'h00; mem['h6D1D]=8'h00; mem['h6D1E]=8'h00; mem['h6D1F]=8'h00;
    mem['h6D20]=8'h00; mem['h6D21]=8'h00; mem['h6D22]=8'h00; mem['h6D23]=8'h00;
    mem['h6D24]=8'h00; mem['h6D25]=8'h00; mem['h6D26]=8'h00; mem['h6D27]=8'h00;
    mem['h6D28]=8'h00; mem['h6D29]=8'h00; mem['h6D2A]=8'h00; mem['h6D2B]=8'h00;
    mem['h6D2C]=8'h00; mem['h6D2D]=8'h00; mem['h6D2E]=8'h00; mem['h6D2F]=8'h00;
    mem['h6D30]=8'h00; mem['h6D31]=8'h00; mem['h6D32]=8'h00; mem['h6D33]=8'h00;
    mem['h6D34]=8'h00; mem['h6D35]=8'h00; mem['h6D36]=8'h00; mem['h6D37]=8'h00;
    mem['h6D38]=8'h00; mem['h6D39]=8'h00; mem['h6D3A]=8'h00; mem['h6D3B]=8'h00;
    mem['h6D3C]=8'h00; mem['h6D3D]=8'h00; mem['h6D3E]=8'h00; mem['h6D3F]=8'h00;
    mem['h6D40]=8'h00; mem['h6D41]=8'h00; mem['h6D42]=8'h00; mem['h6D43]=8'h00;
    mem['h6D44]=8'h00; mem['h6D45]=8'h00; mem['h6D46]=8'h00; mem['h6D47]=8'h00;
    mem['h6D48]=8'h00; mem['h6D49]=8'h00; mem['h6D4A]=8'h00; mem['h6D4B]=8'h00;
    mem['h6D4C]=8'h00; mem['h6D4D]=8'h00; mem['h6D4E]=8'h00; mem['h6D4F]=8'h00;
    mem['h6D50]=8'h00; mem['h6D51]=8'h00; mem['h6D52]=8'h00; mem['h6D53]=8'h00;
    mem['h6D54]=8'h00; mem['h6D55]=8'h00; mem['h6D56]=8'h00; mem['h6D57]=8'h00;
    mem['h6D58]=8'h00; mem['h6D59]=8'h00; mem['h6D5A]=8'h00; mem['h6D5B]=8'h00;
    mem['h6D5C]=8'h00; mem['h6D5D]=8'h00; mem['h6D5E]=8'h00; mem['h6D5F]=8'h00;
    mem['h6D60]=8'h00; mem['h6D61]=8'h00; mem['h6D62]=8'h00; mem['h6D63]=8'h00;
    mem['h6D64]=8'h00; mem['h6D65]=8'h00; mem['h6D66]=8'h00; mem['h6D67]=8'h00;
    mem['h6D68]=8'h00; mem['h6D69]=8'h00; mem['h6D6A]=8'h00; mem['h6D6B]=8'h00;
    mem['h6D6C]=8'h00; mem['h6D6D]=8'h00; mem['h6D6E]=8'h00; mem['h6D6F]=8'h00;
    mem['h6D70]=8'h00; mem['h6D71]=8'h00; mem['h6D72]=8'h00; mem['h6D73]=8'h00;
    mem['h6D74]=8'h00; mem['h6D75]=8'h00; mem['h6D76]=8'h00; mem['h6D77]=8'h00;
    mem['h6D78]=8'h00; mem['h6D79]=8'h00; mem['h6D7A]=8'h00; mem['h6D7B]=8'h00;
    mem['h6D7C]=8'h00; mem['h6D7D]=8'h00; mem['h6D7E]=8'h00; mem['h6D7F]=8'h00;
    mem['h6D80]=8'h00; mem['h6D81]=8'h00; mem['h6D82]=8'h00; mem['h6D83]=8'h00;
    mem['h6D84]=8'h00; mem['h6D85]=8'h00; mem['h6D86]=8'h00; mem['h6D87]=8'h00;
    mem['h6D88]=8'h00; mem['h6D89]=8'h00; mem['h6D8A]=8'h00; mem['h6D8B]=8'h00;
    mem['h6D8C]=8'h00; mem['h6D8D]=8'h00; mem['h6D8E]=8'h00; mem['h6D8F]=8'h00;
    mem['h6D90]=8'h00; mem['h6D91]=8'h00; mem['h6D92]=8'h00; mem['h6D93]=8'h00;
    mem['h6D94]=8'h00; mem['h6D95]=8'h00; mem['h6D96]=8'h00; mem['h6D97]=8'h00;
    mem['h6D98]=8'h00; mem['h6D99]=8'h00; mem['h6D9A]=8'h00; mem['h6D9B]=8'h00;
    mem['h6D9C]=8'h00; mem['h6D9D]=8'h00; mem['h6D9E]=8'h00; mem['h6D9F]=8'h00;
    mem['h6DA0]=8'h00; mem['h6DA1]=8'h00; mem['h6DA2]=8'h00; mem['h6DA3]=8'h00;
    mem['h6DA4]=8'h00; mem['h6DA5]=8'h00; mem['h6DA6]=8'h00; mem['h6DA7]=8'h00;
    mem['h6DA8]=8'h00; mem['h6DA9]=8'h00; mem['h6DAA]=8'h00; mem['h6DAB]=8'h00;
    mem['h6DAC]=8'h00; mem['h6DAD]=8'h00; mem['h6DAE]=8'h00; mem['h6DAF]=8'h00;
    mem['h6DB0]=8'h00; mem['h6DB1]=8'h00; mem['h6DB2]=8'h00; mem['h6DB3]=8'h00;
    mem['h6DB4]=8'h00; mem['h6DB5]=8'h00; mem['h6DB6]=8'h00; mem['h6DB7]=8'h00;
    mem['h6DB8]=8'h00; mem['h6DB9]=8'h00; mem['h6DBA]=8'h00; mem['h6DBB]=8'h00;
    mem['h6DBC]=8'h00; mem['h6DBD]=8'h00; mem['h6DBE]=8'h00; mem['h6DBF]=8'h00;
    mem['h6DC0]=8'h00; mem['h6DC1]=8'h00; mem['h6DC2]=8'h00; mem['h6DC3]=8'h00;
    mem['h6DC4]=8'h00; mem['h6DC5]=8'h00; mem['h6DC6]=8'h00; mem['h6DC7]=8'h00;
    mem['h6DC8]=8'h00; mem['h6DC9]=8'h00; mem['h6DCA]=8'h00; mem['h6DCB]=8'h00;
    mem['h6DCC]=8'h00; mem['h6DCD]=8'h00; mem['h6DCE]=8'h00; mem['h6DCF]=8'h00;
    mem['h6DD0]=8'h00; mem['h6DD1]=8'h00; mem['h6DD2]=8'h00; mem['h6DD3]=8'h00;
    mem['h6DD4]=8'h00; mem['h6DD5]=8'h00; mem['h6DD6]=8'h00; mem['h6DD7]=8'h00;
    mem['h6DD8]=8'h00; mem['h6DD9]=8'h00; mem['h6DDA]=8'h00; mem['h6DDB]=8'h00;
    mem['h6DDC]=8'h00; mem['h6DDD]=8'h00; mem['h6DDE]=8'h00; mem['h6DDF]=8'h00;
    mem['h6DE0]=8'h00; mem['h6DE1]=8'h00; mem['h6DE2]=8'h00; mem['h6DE3]=8'h00;
    mem['h6DE4]=8'h00; mem['h6DE5]=8'h00; mem['h6DE6]=8'h00; mem['h6DE7]=8'h00;
    mem['h6DE8]=8'h00; mem['h6DE9]=8'h00; mem['h6DEA]=8'h00; mem['h6DEB]=8'h00;
    mem['h6DEC]=8'h00; mem['h6DED]=8'h00; mem['h6DEE]=8'h00; mem['h6DEF]=8'h00;
    mem['h6DF0]=8'h00; mem['h6DF1]=8'h00; mem['h6DF2]=8'h00; mem['h6DF3]=8'h00;
    mem['h6DF4]=8'h00; mem['h6DF5]=8'h00; mem['h6DF6]=8'h00; mem['h6DF7]=8'h00;
    mem['h6DF8]=8'h00; mem['h6DF9]=8'h00; mem['h6DFA]=8'h00; mem['h6DFB]=8'h00;
    mem['h6DFC]=8'h00; mem['h6DFD]=8'h00; mem['h6DFE]=8'h00; mem['h6DFF]=8'h00;
    mem['h6E00]=8'h00; mem['h6E01]=8'h00; mem['h6E02]=8'h00; mem['h6E03]=8'h00;
    mem['h6E04]=8'h00; mem['h6E05]=8'h00; mem['h6E06]=8'h00; mem['h6E07]=8'h00;
    mem['h6E08]=8'h00; mem['h6E09]=8'h00; mem['h6E0A]=8'h00; mem['h6E0B]=8'h00;
    mem['h6E0C]=8'h00; mem['h6E0D]=8'h00; mem['h6E0E]=8'h00; mem['h6E0F]=8'h00;
    mem['h6E10]=8'h00; mem['h6E11]=8'h00; mem['h6E12]=8'h00; mem['h6E13]=8'h00;
    mem['h6E14]=8'h00; mem['h6E15]=8'h00; mem['h6E16]=8'h00; mem['h6E17]=8'h00;
    mem['h6E18]=8'h00; mem['h6E19]=8'h00; mem['h6E1A]=8'h00; mem['h6E1B]=8'h00;
    mem['h6E1C]=8'h00; mem['h6E1D]=8'h00; mem['h6E1E]=8'h00; mem['h6E1F]=8'h00;
    mem['h6E20]=8'h00; mem['h6E21]=8'h00; mem['h6E22]=8'h00; mem['h6E23]=8'h00;
    mem['h6E24]=8'h00; mem['h6E25]=8'h00; mem['h6E26]=8'h00; mem['h6E27]=8'h00;
    mem['h6E28]=8'h00; mem['h6E29]=8'h00; mem['h6E2A]=8'h00; mem['h6E2B]=8'h00;
    mem['h6E2C]=8'h00; mem['h6E2D]=8'h00; mem['h6E2E]=8'h00; mem['h6E2F]=8'h00;
    mem['h6E30]=8'h00; mem['h6E31]=8'h00; mem['h6E32]=8'h00; mem['h6E33]=8'h00;
    mem['h6E34]=8'h00; mem['h6E35]=8'h00; mem['h6E36]=8'h00; mem['h6E37]=8'h00;
    mem['h6E38]=8'h00; mem['h6E39]=8'h00; mem['h6E3A]=8'h00; mem['h6E3B]=8'h00;
    mem['h6E3C]=8'h00; mem['h6E3D]=8'h00; mem['h6E3E]=8'h00; mem['h6E3F]=8'h00;
    mem['h6E40]=8'h00; mem['h6E41]=8'h00; mem['h6E42]=8'h00; mem['h6E43]=8'h00;
    mem['h6E44]=8'h00; mem['h6E45]=8'h00; mem['h6E46]=8'h00; mem['h6E47]=8'h00;
    mem['h6E48]=8'h00; mem['h6E49]=8'h00; mem['h6E4A]=8'h00; mem['h6E4B]=8'h00;
    mem['h6E4C]=8'h00; mem['h6E4D]=8'h00; mem['h6E4E]=8'h00; mem['h6E4F]=8'h00;
    mem['h6E50]=8'h00; mem['h6E51]=8'h00; mem['h6E52]=8'h00; mem['h6E53]=8'h00;
    mem['h6E54]=8'h00; mem['h6E55]=8'h00; mem['h6E56]=8'h00; mem['h6E57]=8'h00;
    mem['h6E58]=8'h00; mem['h6E59]=8'h00; mem['h6E5A]=8'h00; mem['h6E5B]=8'h00;
    mem['h6E5C]=8'h00; mem['h6E5D]=8'h00; mem['h6E5E]=8'h00; mem['h6E5F]=8'h00;
    mem['h6E60]=8'h00; mem['h6E61]=8'h00; mem['h6E62]=8'h00; mem['h6E63]=8'h00;
    mem['h6E64]=8'h00; mem['h6E65]=8'h00; mem['h6E66]=8'h00; mem['h6E67]=8'h00;
    mem['h6E68]=8'h00; mem['h6E69]=8'h00; mem['h6E6A]=8'h00; mem['h6E6B]=8'h00;
    mem['h6E6C]=8'h00; mem['h6E6D]=8'h00; mem['h6E6E]=8'h00; mem['h6E6F]=8'h00;
    mem['h6E70]=8'h00; mem['h6E71]=8'h00; mem['h6E72]=8'h00; mem['h6E73]=8'h00;
    mem['h6E74]=8'h00; mem['h6E75]=8'h00; mem['h6E76]=8'h00; mem['h6E77]=8'h00;
    mem['h6E78]=8'h00; mem['h6E79]=8'h00; mem['h6E7A]=8'h00; mem['h6E7B]=8'h00;
    mem['h6E7C]=8'h00; mem['h6E7D]=8'h00; mem['h6E7E]=8'h00; mem['h6E7F]=8'h00;
    mem['h6E80]=8'h00; mem['h6E81]=8'h00; mem['h6E82]=8'h00; mem['h6E83]=8'h00;
    mem['h6E84]=8'h00; mem['h6E85]=8'h00; mem['h6E86]=8'h00; mem['h6E87]=8'h00;
    mem['h6E88]=8'h00; mem['h6E89]=8'h00; mem['h6E8A]=8'h00; mem['h6E8B]=8'h00;
    mem['h6E8C]=8'h00; mem['h6E8D]=8'h00; mem['h6E8E]=8'h00; mem['h6E8F]=8'h00;
    mem['h6E90]=8'h00; mem['h6E91]=8'h00; mem['h6E92]=8'h00; mem['h6E93]=8'h00;
    mem['h6E94]=8'h00; mem['h6E95]=8'h00; mem['h6E96]=8'h00; mem['h6E97]=8'h00;
    mem['h6E98]=8'h00; mem['h6E99]=8'h00; mem['h6E9A]=8'h00; mem['h6E9B]=8'h00;
    mem['h6E9C]=8'h00; mem['h6E9D]=8'h00; mem['h6E9E]=8'h00; mem['h6E9F]=8'h00;
    mem['h6EA0]=8'h00; mem['h6EA1]=8'h00; mem['h6EA2]=8'h00; mem['h6EA3]=8'h00;
    mem['h6EA4]=8'h00; mem['h6EA5]=8'h00; mem['h6EA6]=8'h00; mem['h6EA7]=8'h00;
    mem['h6EA8]=8'h00; mem['h6EA9]=8'h00; mem['h6EAA]=8'h00; mem['h6EAB]=8'h00;
    mem['h6EAC]=8'h00; mem['h6EAD]=8'h00; mem['h6EAE]=8'h00; mem['h6EAF]=8'h00;
    mem['h6EB0]=8'h00; mem['h6EB1]=8'h00; mem['h6EB2]=8'h00; mem['h6EB3]=8'h00;
    mem['h6EB4]=8'h00; mem['h6EB5]=8'h00; mem['h6EB6]=8'h00; mem['h6EB7]=8'h00;
    mem['h6EB8]=8'h00; mem['h6EB9]=8'h00; mem['h6EBA]=8'h00; mem['h6EBB]=8'h00;
    mem['h6EBC]=8'h00; mem['h6EBD]=8'h00; mem['h6EBE]=8'h00; mem['h6EBF]=8'h00;
    mem['h6EC0]=8'h00; mem['h6EC1]=8'h00; mem['h6EC2]=8'h00; mem['h6EC3]=8'h00;
    mem['h6EC4]=8'h00; mem['h6EC5]=8'h00; mem['h6EC6]=8'h00; mem['h6EC7]=8'h00;
    mem['h6EC8]=8'h00; mem['h6EC9]=8'h00; mem['h6ECA]=8'h00; mem['h6ECB]=8'h00;
    mem['h6ECC]=8'h00; mem['h6ECD]=8'h00; mem['h6ECE]=8'h00; mem['h6ECF]=8'h00;
    mem['h6ED0]=8'h00; mem['h6ED1]=8'h00; mem['h6ED2]=8'h00; mem['h6ED3]=8'h00;
    mem['h6ED4]=8'h00; mem['h6ED5]=8'h00; mem['h6ED6]=8'h00; mem['h6ED7]=8'h00;
    mem['h6ED8]=8'h00; mem['h6ED9]=8'h00; mem['h6EDA]=8'h00; mem['h6EDB]=8'h00;
    mem['h6EDC]=8'h00; mem['h6EDD]=8'h00; mem['h6EDE]=8'h00; mem['h6EDF]=8'h00;
    mem['h6EE0]=8'h00; mem['h6EE1]=8'h00; mem['h6EE2]=8'h00; mem['h6EE3]=8'h00;
    mem['h6EE4]=8'h00; mem['h6EE5]=8'h00; mem['h6EE6]=8'h00; mem['h6EE7]=8'h00;
    mem['h6EE8]=8'h00; mem['h6EE9]=8'h00; mem['h6EEA]=8'h00; mem['h6EEB]=8'h00;
    mem['h6EEC]=8'h00; mem['h6EED]=8'h00; mem['h6EEE]=8'h00; mem['h6EEF]=8'h00;
    mem['h6EF0]=8'h00; mem['h6EF1]=8'h00; mem['h6EF2]=8'h00; mem['h6EF3]=8'h00;
    mem['h6EF4]=8'h00; mem['h6EF5]=8'h00; mem['h6EF6]=8'h00; mem['h6EF7]=8'h00;
    mem['h6EF8]=8'h00; mem['h6EF9]=8'h00; mem['h6EFA]=8'h00; mem['h6EFB]=8'h00;
    mem['h6EFC]=8'h00; mem['h6EFD]=8'h00; mem['h6EFE]=8'h00; mem['h6EFF]=8'h00;
    mem['h6F00]=8'h00; mem['h6F01]=8'h00; mem['h6F02]=8'h00; mem['h6F03]=8'h00;
    mem['h6F04]=8'h00; mem['h6F05]=8'h00; mem['h6F06]=8'h00; mem['h6F07]=8'h00;
    mem['h6F08]=8'h00; mem['h6F09]=8'h00; mem['h6F0A]=8'h00; mem['h6F0B]=8'h00;
    mem['h6F0C]=8'h00; mem['h6F0D]=8'h00; mem['h6F0E]=8'h00; mem['h6F0F]=8'h00;
    mem['h6F10]=8'h00; mem['h6F11]=8'h00; mem['h6F12]=8'h00; mem['h6F13]=8'h00;
    mem['h6F14]=8'h00; mem['h6F15]=8'h00; mem['h6F16]=8'h00; mem['h6F17]=8'h00;
    mem['h6F18]=8'h00; mem['h6F19]=8'h00; mem['h6F1A]=8'h00; mem['h6F1B]=8'h00;
    mem['h6F1C]=8'h00; mem['h6F1D]=8'h00; mem['h6F1E]=8'h00; mem['h6F1F]=8'h00;
    mem['h6F20]=8'h00; mem['h6F21]=8'h00; mem['h6F22]=8'h00; mem['h6F23]=8'h00;
    mem['h6F24]=8'h00; mem['h6F25]=8'h00; mem['h6F26]=8'h00; mem['h6F27]=8'h00;
    mem['h6F28]=8'h00; mem['h6F29]=8'h00; mem['h6F2A]=8'h00; mem['h6F2B]=8'h00;
    mem['h6F2C]=8'h00; mem['h6F2D]=8'h00; mem['h6F2E]=8'h00; mem['h6F2F]=8'h00;
    mem['h6F30]=8'h00; mem['h6F31]=8'h00; mem['h6F32]=8'h00; mem['h6F33]=8'h00;
    mem['h6F34]=8'h00; mem['h6F35]=8'h00; mem['h6F36]=8'h00; mem['h6F37]=8'h00;
    mem['h6F38]=8'h00; mem['h6F39]=8'h00; mem['h6F3A]=8'h00; mem['h6F3B]=8'h00;
    mem['h6F3C]=8'h00; mem['h6F3D]=8'h00; mem['h6F3E]=8'h00; mem['h6F3F]=8'h00;
    mem['h6F40]=8'h00; mem['h6F41]=8'h00; mem['h6F42]=8'h00; mem['h6F43]=8'h00;
    mem['h6F44]=8'h00; mem['h6F45]=8'h00; mem['h6F46]=8'h00; mem['h6F47]=8'h00;
    mem['h6F48]=8'h00; mem['h6F49]=8'h00; mem['h6F4A]=8'h00; mem['h6F4B]=8'h00;
    mem['h6F4C]=8'h00; mem['h6F4D]=8'h00; mem['h6F4E]=8'h00; mem['h6F4F]=8'h00;
    mem['h6F50]=8'h00; mem['h6F51]=8'h00; mem['h6F52]=8'h00; mem['h6F53]=8'h00;
    mem['h6F54]=8'h00; mem['h6F55]=8'h00; mem['h6F56]=8'h00; mem['h6F57]=8'h00;
    mem['h6F58]=8'h00; mem['h6F59]=8'h00; mem['h6F5A]=8'h00; mem['h6F5B]=8'h00;
    mem['h6F5C]=8'h00; mem['h6F5D]=8'h00; mem['h6F5E]=8'h00; mem['h6F5F]=8'h00;
    mem['h6F60]=8'h00; mem['h6F61]=8'h00; mem['h6F62]=8'h00; mem['h6F63]=8'h00;
    mem['h6F64]=8'h00; mem['h6F65]=8'h00; mem['h6F66]=8'h00; mem['h6F67]=8'h00;
    mem['h6F68]=8'h00; mem['h6F69]=8'h00; mem['h6F6A]=8'h00; mem['h6F6B]=8'h00;
    mem['h6F6C]=8'h00; mem['h6F6D]=8'h00; mem['h6F6E]=8'h00; mem['h6F6F]=8'h00;
    mem['h6F70]=8'h00; mem['h6F71]=8'h00; mem['h6F72]=8'h00; mem['h6F73]=8'h00;
    mem['h6F74]=8'h00; mem['h6F75]=8'h00; mem['h6F76]=8'h00; mem['h6F77]=8'h00;
    mem['h6F78]=8'h00; mem['h6F79]=8'h00; mem['h6F7A]=8'h00; mem['h6F7B]=8'h00;
    mem['h6F7C]=8'h00; mem['h6F7D]=8'h00; mem['h6F7E]=8'h00; mem['h6F7F]=8'h00;
    mem['h6F80]=8'h00; mem['h6F81]=8'h00; mem['h6F82]=8'h00; mem['h6F83]=8'h00;
    mem['h6F84]=8'h00; mem['h6F85]=8'h00; mem['h6F86]=8'h00; mem['h6F87]=8'h00;
    mem['h6F88]=8'h00; mem['h6F89]=8'h00; mem['h6F8A]=8'h00; mem['h6F8B]=8'h00;
    mem['h6F8C]=8'h00; mem['h6F8D]=8'h00; mem['h6F8E]=8'h00; mem['h6F8F]=8'h00;
    mem['h6F90]=8'h00; mem['h6F91]=8'h00; mem['h6F92]=8'h00; mem['h6F93]=8'h00;
    mem['h6F94]=8'h00; mem['h6F95]=8'h00; mem['h6F96]=8'h00; mem['h6F97]=8'h00;
    mem['h6F98]=8'h00; mem['h6F99]=8'h00; mem['h6F9A]=8'h00; mem['h6F9B]=8'h00;
    mem['h6F9C]=8'h00; mem['h6F9D]=8'h00; mem['h6F9E]=8'h00; mem['h6F9F]=8'h00;
    mem['h6FA0]=8'h00; mem['h6FA1]=8'h00; mem['h6FA2]=8'h00; mem['h6FA3]=8'h00;
    mem['h6FA4]=8'h00; mem['h6FA5]=8'h00; mem['h6FA6]=8'h00; mem['h6FA7]=8'h00;
    mem['h6FA8]=8'h00; mem['h6FA9]=8'h00; mem['h6FAA]=8'h00; mem['h6FAB]=8'h00;
    mem['h6FAC]=8'h00; mem['h6FAD]=8'h00; mem['h6FAE]=8'h00; mem['h6FAF]=8'h00;
    mem['h6FB0]=8'h00; mem['h6FB1]=8'h00; mem['h6FB2]=8'h00; mem['h6FB3]=8'h00;
    mem['h6FB4]=8'h00; mem['h6FB5]=8'h00; mem['h6FB6]=8'h00; mem['h6FB7]=8'h00;
    mem['h6FB8]=8'h00; mem['h6FB9]=8'h00; mem['h6FBA]=8'h00; mem['h6FBB]=8'h00;
    mem['h6FBC]=8'h00; mem['h6FBD]=8'h00; mem['h6FBE]=8'h00; mem['h6FBF]=8'h00;
    mem['h6FC0]=8'h00; mem['h6FC1]=8'h00; mem['h6FC2]=8'h00; mem['h6FC3]=8'h00;
    mem['h6FC4]=8'h00; mem['h6FC5]=8'h00; mem['h6FC6]=8'h00; mem['h6FC7]=8'h00;
    mem['h6FC8]=8'h00; mem['h6FC9]=8'h00; mem['h6FCA]=8'h00; mem['h6FCB]=8'h00;
    mem['h6FCC]=8'h00; mem['h6FCD]=8'h00; mem['h6FCE]=8'h00; mem['h6FCF]=8'h00;
    mem['h6FD0]=8'h00; mem['h6FD1]=8'h00; mem['h6FD2]=8'h00; mem['h6FD3]=8'h00;
    mem['h6FD4]=8'h00; mem['h6FD5]=8'h00; mem['h6FD6]=8'h00; mem['h6FD7]=8'h00;
    mem['h6FD8]=8'h00; mem['h6FD9]=8'h00; mem['h6FDA]=8'h00; mem['h6FDB]=8'h00;
    mem['h6FDC]=8'h00; mem['h6FDD]=8'h00; mem['h6FDE]=8'h00; mem['h6FDF]=8'h00;
    mem['h6FE0]=8'h00; mem['h6FE1]=8'h00; mem['h6FE2]=8'h00; mem['h6FE3]=8'h00;
    mem['h6FE4]=8'h00; mem['h6FE5]=8'h00; mem['h6FE6]=8'h00; mem['h6FE7]=8'h00;
    mem['h6FE8]=8'h00; mem['h6FE9]=8'h00; mem['h6FEA]=8'h00; mem['h6FEB]=8'h00;
    mem['h6FEC]=8'h00; mem['h6FED]=8'h00; mem['h6FEE]=8'h00; mem['h6FEF]=8'h00;
    mem['h6FF0]=8'h00; mem['h6FF1]=8'h00; mem['h6FF2]=8'h00; mem['h6FF3]=8'h00;
    mem['h6FF4]=8'h00; mem['h6FF5]=8'h00; mem['h6FF6]=8'h00; mem['h6FF7]=8'h00;
    mem['h6FF8]=8'h00; mem['h6FF9]=8'h00; mem['h6FFA]=8'h00; mem['h6FFB]=8'h00;
    mem['h6FFC]=8'h00; mem['h6FFD]=8'h00; mem['h6FFE]=8'h00; mem['h6FFF]=8'h00;
    mem['h7000]=8'h00; mem['h7001]=8'h00; mem['h7002]=8'h00; mem['h7003]=8'h00;
    mem['h7004]=8'h00; mem['h7005]=8'h00; mem['h7006]=8'h00; mem['h7007]=8'h00;
    mem['h7008]=8'h00; mem['h7009]=8'h00; mem['h700A]=8'h00; mem['h700B]=8'h00;
    mem['h700C]=8'h00; mem['h700D]=8'h00; mem['h700E]=8'h00; mem['h700F]=8'h00;
    mem['h7010]=8'h00; mem['h7011]=8'h00; mem['h7012]=8'h00; mem['h7013]=8'h00;
    mem['h7014]=8'h00; mem['h7015]=8'h00; mem['h7016]=8'h00; mem['h7017]=8'h00;
    mem['h7018]=8'h00; mem['h7019]=8'h00; mem['h701A]=8'h00; mem['h701B]=8'h00;
    mem['h701C]=8'h00; mem['h701D]=8'h00; mem['h701E]=8'h00; mem['h701F]=8'h00;
    mem['h7020]=8'h00; mem['h7021]=8'h00; mem['h7022]=8'h00; mem['h7023]=8'h00;
    mem['h7024]=8'h00; mem['h7025]=8'h00; mem['h7026]=8'h00; mem['h7027]=8'h00;
    mem['h7028]=8'h00; mem['h7029]=8'h00; mem['h702A]=8'h00; mem['h702B]=8'h00;
    mem['h702C]=8'h00; mem['h702D]=8'h00; mem['h702E]=8'h00; mem['h702F]=8'h00;
    mem['h7030]=8'h00; mem['h7031]=8'h00; mem['h7032]=8'h00; mem['h7033]=8'h00;
    mem['h7034]=8'h00; mem['h7035]=8'h00; mem['h7036]=8'h00; mem['h7037]=8'h00;
    mem['h7038]=8'h00; mem['h7039]=8'h00; mem['h703A]=8'h00; mem['h703B]=8'h00;
    mem['h703C]=8'h00; mem['h703D]=8'h00; mem['h703E]=8'h00; mem['h703F]=8'h00;
    mem['h7040]=8'h00; mem['h7041]=8'h00; mem['h7042]=8'h00; mem['h7043]=8'h00;
    mem['h7044]=8'h00; mem['h7045]=8'h00; mem['h7046]=8'h00; mem['h7047]=8'h00;
    mem['h7048]=8'h00; mem['h7049]=8'h00; mem['h704A]=8'h00; mem['h704B]=8'h00;
    mem['h704C]=8'h00; mem['h704D]=8'h00; mem['h704E]=8'h00; mem['h704F]=8'h00;
    mem['h7050]=8'h00; mem['h7051]=8'h00; mem['h7052]=8'h00; mem['h7053]=8'h00;
    mem['h7054]=8'h00; mem['h7055]=8'h00; mem['h7056]=8'h00; mem['h7057]=8'h00;
    mem['h7058]=8'h00; mem['h7059]=8'h00; mem['h705A]=8'h00; mem['h705B]=8'h00;
    mem['h705C]=8'h00; mem['h705D]=8'h00; mem['h705E]=8'h00; mem['h705F]=8'h00;
    mem['h7060]=8'h00; mem['h7061]=8'h00; mem['h7062]=8'h00; mem['h7063]=8'h00;
    mem['h7064]=8'h00; mem['h7065]=8'h00; mem['h7066]=8'h00; mem['h7067]=8'h00;
    mem['h7068]=8'h00; mem['h7069]=8'h00; mem['h706A]=8'h00; mem['h706B]=8'h00;
    mem['h706C]=8'h00; mem['h706D]=8'h00; mem['h706E]=8'h00; mem['h706F]=8'h00;
    mem['h7070]=8'h00; mem['h7071]=8'h00; mem['h7072]=8'h00; mem['h7073]=8'h00;
    mem['h7074]=8'h00; mem['h7075]=8'h00; mem['h7076]=8'h00; mem['h7077]=8'h00;
    mem['h7078]=8'h00; mem['h7079]=8'h00; mem['h707A]=8'h00; mem['h707B]=8'h00;
    mem['h707C]=8'h00; mem['h707D]=8'h00; mem['h707E]=8'h00; mem['h707F]=8'h00;
    mem['h7080]=8'h00; mem['h7081]=8'h00; mem['h7082]=8'h00; mem['h7083]=8'h00;
    mem['h7084]=8'h00; mem['h7085]=8'h00; mem['h7086]=8'h00; mem['h7087]=8'h00;
    mem['h7088]=8'h00; mem['h7089]=8'h00; mem['h708A]=8'h00; mem['h708B]=8'h00;
    mem['h708C]=8'h00; mem['h708D]=8'h00; mem['h708E]=8'h00; mem['h708F]=8'h00;
    mem['h7090]=8'h00; mem['h7091]=8'h00; mem['h7092]=8'h00; mem['h7093]=8'h00;
    mem['h7094]=8'h00; mem['h7095]=8'h00; mem['h7096]=8'h00; mem['h7097]=8'h00;
    mem['h7098]=8'h00; mem['h7099]=8'h00; mem['h709A]=8'h00; mem['h709B]=8'h00;
    mem['h709C]=8'h00; mem['h709D]=8'h00; mem['h709E]=8'h00; mem['h709F]=8'h00;
    mem['h70A0]=8'h00; mem['h70A1]=8'h00; mem['h70A2]=8'h00; mem['h70A3]=8'h00;
    mem['h70A4]=8'h00; mem['h70A5]=8'h00; mem['h70A6]=8'h00; mem['h70A7]=8'h00;
    mem['h70A8]=8'h00; mem['h70A9]=8'h00; mem['h70AA]=8'h00; mem['h70AB]=8'h00;
    mem['h70AC]=8'h00; mem['h70AD]=8'h00; mem['h70AE]=8'h00; mem['h70AF]=8'h00;
    mem['h70B0]=8'h00; mem['h70B1]=8'h00; mem['h70B2]=8'h00; mem['h70B3]=8'h00;
    mem['h70B4]=8'h00; mem['h70B5]=8'h00; mem['h70B6]=8'h00; mem['h70B7]=8'h00;
    mem['h70B8]=8'h00; mem['h70B9]=8'h00; mem['h70BA]=8'h00; mem['h70BB]=8'h00;
    mem['h70BC]=8'h00; mem['h70BD]=8'h00; mem['h70BE]=8'h00; mem['h70BF]=8'h00;
    mem['h70C0]=8'h00; mem['h70C1]=8'h00; mem['h70C2]=8'h00; mem['h70C3]=8'h00;
    mem['h70C4]=8'h00; mem['h70C5]=8'h00; mem['h70C6]=8'h00; mem['h70C7]=8'h00;
    mem['h70C8]=8'h00; mem['h70C9]=8'h00; mem['h70CA]=8'h00; mem['h70CB]=8'h00;
    mem['h70CC]=8'h00; mem['h70CD]=8'h00; mem['h70CE]=8'h00; mem['h70CF]=8'h00;
    mem['h70D0]=8'h00; mem['h70D1]=8'h00; mem['h70D2]=8'h00; mem['h70D3]=8'h00;
    mem['h70D4]=8'h00; mem['h70D5]=8'h00; mem['h70D6]=8'h00; mem['h70D7]=8'h00;
    mem['h70D8]=8'h00; mem['h70D9]=8'h00; mem['h70DA]=8'h00; mem['h70DB]=8'h00;
    mem['h70DC]=8'h00; mem['h70DD]=8'h00; mem['h70DE]=8'h00; mem['h70DF]=8'h00;
    mem['h70E0]=8'h00; mem['h70E1]=8'h00; mem['h70E2]=8'h00; mem['h70E3]=8'h00;
    mem['h70E4]=8'h00; mem['h70E5]=8'h00; mem['h70E6]=8'h00; mem['h70E7]=8'h00;
    mem['h70E8]=8'h00; mem['h70E9]=8'h00; mem['h70EA]=8'h00; mem['h70EB]=8'h00;
    mem['h70EC]=8'h00; mem['h70ED]=8'h00; mem['h70EE]=8'h00; mem['h70EF]=8'h00;
    mem['h70F0]=8'h00; mem['h70F1]=8'h00; mem['h70F2]=8'h00; mem['h70F3]=8'h00;
    mem['h70F4]=8'h00; mem['h70F5]=8'h00; mem['h70F6]=8'h00; mem['h70F7]=8'h00;
    mem['h70F8]=8'h00; mem['h70F9]=8'h00; mem['h70FA]=8'h00; mem['h70FB]=8'h00;
    mem['h70FC]=8'h00; mem['h70FD]=8'h00; mem['h70FE]=8'h00; mem['h70FF]=8'h00;
    mem['h7100]=8'h00; mem['h7101]=8'h00; mem['h7102]=8'h00; mem['h7103]=8'h00;
    mem['h7104]=8'h00; mem['h7105]=8'h00; mem['h7106]=8'h00; mem['h7107]=8'h00;
    mem['h7108]=8'h00; mem['h7109]=8'h00; mem['h710A]=8'h00; mem['h710B]=8'h00;
    mem['h710C]=8'h00; mem['h710D]=8'h00; mem['h710E]=8'h00; mem['h710F]=8'h00;
    mem['h7110]=8'h00; mem['h7111]=8'h00; mem['h7112]=8'h00; mem['h7113]=8'h00;
    mem['h7114]=8'h00; mem['h7115]=8'h00; mem['h7116]=8'h00; mem['h7117]=8'h00;
    mem['h7118]=8'h00; mem['h7119]=8'h00; mem['h711A]=8'h00; mem['h711B]=8'h00;
    mem['h711C]=8'h00; mem['h711D]=8'h00; mem['h711E]=8'h00; mem['h711F]=8'h00;
    mem['h7120]=8'h00; mem['h7121]=8'h00; mem['h7122]=8'h00; mem['h7123]=8'h00;
    mem['h7124]=8'h00; mem['h7125]=8'h00; mem['h7126]=8'h00; mem['h7127]=8'h00;
    mem['h7128]=8'h00; mem['h7129]=8'h00; mem['h712A]=8'h00; mem['h712B]=8'h00;
    mem['h712C]=8'h00; mem['h712D]=8'h00; mem['h712E]=8'h00; mem['h712F]=8'h00;
    mem['h7130]=8'h00; mem['h7131]=8'h00; mem['h7132]=8'h00; mem['h7133]=8'h00;
    mem['h7134]=8'h00; mem['h7135]=8'h00; mem['h7136]=8'h00; mem['h7137]=8'h00;
    mem['h7138]=8'h00; mem['h7139]=8'h00; mem['h713A]=8'h00; mem['h713B]=8'h00;
    mem['h713C]=8'h00; mem['h713D]=8'h00; mem['h713E]=8'h00; mem['h713F]=8'h00;
    mem['h7140]=8'h00; mem['h7141]=8'h00; mem['h7142]=8'h00; mem['h7143]=8'h00;
    mem['h7144]=8'h00; mem['h7145]=8'h00; mem['h7146]=8'h00; mem['h7147]=8'h00;
    mem['h7148]=8'h00; mem['h7149]=8'h00; mem['h714A]=8'h00; mem['h714B]=8'h00;
    mem['h714C]=8'h00; mem['h714D]=8'h00; mem['h714E]=8'h00; mem['h714F]=8'h00;
    mem['h7150]=8'h00; mem['h7151]=8'h00; mem['h7152]=8'h00; mem['h7153]=8'h00;
    mem['h7154]=8'h00; mem['h7155]=8'h00; mem['h7156]=8'h00; mem['h7157]=8'h00;
    mem['h7158]=8'h00; mem['h7159]=8'h00; mem['h715A]=8'h00; mem['h715B]=8'h00;
    mem['h715C]=8'h00; mem['h715D]=8'h00; mem['h715E]=8'h00; mem['h715F]=8'h00;
    mem['h7160]=8'h00; mem['h7161]=8'h00; mem['h7162]=8'h00; mem['h7163]=8'h00;
    mem['h7164]=8'h00; mem['h7165]=8'h00; mem['h7166]=8'h00; mem['h7167]=8'h00;
    mem['h7168]=8'h00; mem['h7169]=8'h00; mem['h716A]=8'h00; mem['h716B]=8'h00;
    mem['h716C]=8'h00; mem['h716D]=8'h00; mem['h716E]=8'h00; mem['h716F]=8'h00;
    mem['h7170]=8'h00; mem['h7171]=8'h00; mem['h7172]=8'h00; mem['h7173]=8'h00;
    mem['h7174]=8'h00; mem['h7175]=8'h00; mem['h7176]=8'h00; mem['h7177]=8'h00;
    mem['h7178]=8'h00; mem['h7179]=8'h00; mem['h717A]=8'h00; mem['h717B]=8'h00;
    mem['h717C]=8'h00; mem['h717D]=8'h00; mem['h717E]=8'h00; mem['h717F]=8'h00;
    mem['h7180]=8'h00; mem['h7181]=8'h00; mem['h7182]=8'h00; mem['h7183]=8'h00;
    mem['h7184]=8'h00; mem['h7185]=8'h00; mem['h7186]=8'h00; mem['h7187]=8'h00;
    mem['h7188]=8'h00; mem['h7189]=8'h00; mem['h718A]=8'h00; mem['h718B]=8'h00;
    mem['h718C]=8'h00; mem['h718D]=8'h00; mem['h718E]=8'h00; mem['h718F]=8'h00;
    mem['h7190]=8'h00; mem['h7191]=8'h00; mem['h7192]=8'h00; mem['h7193]=8'h00;
    mem['h7194]=8'h00; mem['h7195]=8'h00; mem['h7196]=8'h00; mem['h7197]=8'h00;
    mem['h7198]=8'h00; mem['h7199]=8'h00; mem['h719A]=8'h00; mem['h719B]=8'h00;
    mem['h719C]=8'h00; mem['h719D]=8'h00; mem['h719E]=8'h00; mem['h719F]=8'h00;
    mem['h71A0]=8'h00; mem['h71A1]=8'h00; mem['h71A2]=8'h00; mem['h71A3]=8'h00;
    mem['h71A4]=8'h00; mem['h71A5]=8'h00; mem['h71A6]=8'h00; mem['h71A7]=8'h00;
    mem['h71A8]=8'h00; mem['h71A9]=8'h00; mem['h71AA]=8'h00; mem['h71AB]=8'h00;
    mem['h71AC]=8'h00; mem['h71AD]=8'h00; mem['h71AE]=8'h00; mem['h71AF]=8'h00;
    mem['h71B0]=8'h00; mem['h71B1]=8'h00; mem['h71B2]=8'h00; mem['h71B3]=8'h00;
    mem['h71B4]=8'h00; mem['h71B5]=8'h00; mem['h71B6]=8'h00; mem['h71B7]=8'h00;
    mem['h71B8]=8'h00; mem['h71B9]=8'h00; mem['h71BA]=8'h00; mem['h71BB]=8'h00;
    mem['h71BC]=8'h00; mem['h71BD]=8'h00; mem['h71BE]=8'h00; mem['h71BF]=8'h00;
    mem['h71C0]=8'h00; mem['h71C1]=8'h00; mem['h71C2]=8'h00; mem['h71C3]=8'h00;
    mem['h71C4]=8'h00; mem['h71C5]=8'h00; mem['h71C6]=8'h00; mem['h71C7]=8'h00;
    mem['h71C8]=8'h00; mem['h71C9]=8'h00; mem['h71CA]=8'h00; mem['h71CB]=8'h00;
    mem['h71CC]=8'h00; mem['h71CD]=8'h00; mem['h71CE]=8'h00; mem['h71CF]=8'h00;
    mem['h71D0]=8'h00; mem['h71D1]=8'h00; mem['h71D2]=8'h00; mem['h71D3]=8'h00;
    mem['h71D4]=8'h00; mem['h71D5]=8'h00; mem['h71D6]=8'h00; mem['h71D7]=8'h00;
    mem['h71D8]=8'h00; mem['h71D9]=8'h00; mem['h71DA]=8'h00; mem['h71DB]=8'h00;
    mem['h71DC]=8'h00; mem['h71DD]=8'h00; mem['h71DE]=8'h00; mem['h71DF]=8'h00;
    mem['h71E0]=8'h00; mem['h71E1]=8'h00; mem['h71E2]=8'h00; mem['h71E3]=8'h00;
    mem['h71E4]=8'h00; mem['h71E5]=8'h00; mem['h71E6]=8'h00; mem['h71E7]=8'h00;
    mem['h71E8]=8'h00; mem['h71E9]=8'h00; mem['h71EA]=8'h00; mem['h71EB]=8'h00;
    mem['h71EC]=8'h00; mem['h71ED]=8'h00; mem['h71EE]=8'h00; mem['h71EF]=8'h00;
    mem['h71F0]=8'h00; mem['h71F1]=8'h00; mem['h71F2]=8'h00; mem['h71F3]=8'h00;
    mem['h71F4]=8'h00; mem['h71F5]=8'h00; mem['h71F6]=8'h00; mem['h71F7]=8'h00;
    mem['h71F8]=8'h00; mem['h71F9]=8'h00; mem['h71FA]=8'h00; mem['h71FB]=8'h00;
    mem['h71FC]=8'h00; mem['h71FD]=8'h00; mem['h71FE]=8'h00; mem['h71FF]=8'h00;
    mem['h7200]=8'h00; mem['h7201]=8'h00; mem['h7202]=8'h00; mem['h7203]=8'h00;
    mem['h7204]=8'h00; mem['h7205]=8'h00; mem['h7206]=8'h00; mem['h7207]=8'h00;
    mem['h7208]=8'h00; mem['h7209]=8'h00; mem['h720A]=8'h00; mem['h720B]=8'h00;
    mem['h720C]=8'h00; mem['h720D]=8'h00; mem['h720E]=8'h00; mem['h720F]=8'h00;
    mem['h7210]=8'h00; mem['h7211]=8'h00; mem['h7212]=8'h00; mem['h7213]=8'h00;
    mem['h7214]=8'h00; mem['h7215]=8'h00; mem['h7216]=8'h00; mem['h7217]=8'h00;
    mem['h7218]=8'h00; mem['h7219]=8'h00; mem['h721A]=8'h00; mem['h721B]=8'h00;
    mem['h721C]=8'h00; mem['h721D]=8'h00; mem['h721E]=8'h00; mem['h721F]=8'h00;
    mem['h7220]=8'h00; mem['h7221]=8'h00; mem['h7222]=8'h00; mem['h7223]=8'h00;
    mem['h7224]=8'h00; mem['h7225]=8'h00; mem['h7226]=8'h00; mem['h7227]=8'h00;
    mem['h7228]=8'h00; mem['h7229]=8'h00; mem['h722A]=8'h00; mem['h722B]=8'h00;
    mem['h722C]=8'h00; mem['h722D]=8'h00; mem['h722E]=8'h00; mem['h722F]=8'h00;
    mem['h7230]=8'h00; mem['h7231]=8'h00; mem['h7232]=8'h00; mem['h7233]=8'h00;
    mem['h7234]=8'h00; mem['h7235]=8'h00; mem['h7236]=8'h00; mem['h7237]=8'h00;
    mem['h7238]=8'h00; mem['h7239]=8'h00; mem['h723A]=8'h00; mem['h723B]=8'h00;
    mem['h723C]=8'h00; mem['h723D]=8'h00; mem['h723E]=8'h00; mem['h723F]=8'h00;
    mem['h7240]=8'h00; mem['h7241]=8'h00; mem['h7242]=8'h00; mem['h7243]=8'h00;
    mem['h7244]=8'h00; mem['h7245]=8'h00; mem['h7246]=8'h00; mem['h7247]=8'h00;
    mem['h7248]=8'h00; mem['h7249]=8'h00; mem['h724A]=8'h00; mem['h724B]=8'h00;
    mem['h724C]=8'h00; mem['h724D]=8'h00; mem['h724E]=8'h00; mem['h724F]=8'h00;
    mem['h7250]=8'h00; mem['h7251]=8'h00; mem['h7252]=8'h00; mem['h7253]=8'h00;
    mem['h7254]=8'h00; mem['h7255]=8'h00; mem['h7256]=8'h00; mem['h7257]=8'h00;
    mem['h7258]=8'h00; mem['h7259]=8'h00; mem['h725A]=8'h00; mem['h725B]=8'h00;
    mem['h725C]=8'h00; mem['h725D]=8'h00; mem['h725E]=8'h00; mem['h725F]=8'h00;
    mem['h7260]=8'h00; mem['h7261]=8'h00; mem['h7262]=8'h00; mem['h7263]=8'h00;
    mem['h7264]=8'h00; mem['h7265]=8'h00; mem['h7266]=8'h00; mem['h7267]=8'h00;
    mem['h7268]=8'h00; mem['h7269]=8'h00; mem['h726A]=8'h00; mem['h726B]=8'h00;
    mem['h726C]=8'h00; mem['h726D]=8'h00; mem['h726E]=8'h00; mem['h726F]=8'h00;
    mem['h7270]=8'h00; mem['h7271]=8'h00; mem['h7272]=8'h00; mem['h7273]=8'h00;
    mem['h7274]=8'h00; mem['h7275]=8'h00; mem['h7276]=8'h00; mem['h7277]=8'h00;
    mem['h7278]=8'h00; mem['h7279]=8'h00; mem['h727A]=8'h00; mem['h727B]=8'h00;
    mem['h727C]=8'h00; mem['h727D]=8'h00; mem['h727E]=8'h00; mem['h727F]=8'h00;
    mem['h7280]=8'h00; mem['h7281]=8'h00; mem['h7282]=8'h00; mem['h7283]=8'h00;
    mem['h7284]=8'h00; mem['h7285]=8'h00; mem['h7286]=8'h00; mem['h7287]=8'h00;
    mem['h7288]=8'h00; mem['h7289]=8'h00; mem['h728A]=8'h00; mem['h728B]=8'h00;
    mem['h728C]=8'h00; mem['h728D]=8'h00; mem['h728E]=8'h00; mem['h728F]=8'h00;
    mem['h7290]=8'h00; mem['h7291]=8'h00; mem['h7292]=8'h00; mem['h7293]=8'h00;
    mem['h7294]=8'h00; mem['h7295]=8'h00; mem['h7296]=8'h00; mem['h7297]=8'h00;
    mem['h7298]=8'h00; mem['h7299]=8'h00; mem['h729A]=8'h00; mem['h729B]=8'h00;
    mem['h729C]=8'h00; mem['h729D]=8'h00; mem['h729E]=8'h00; mem['h729F]=8'h00;
    mem['h72A0]=8'h00; mem['h72A1]=8'h00; mem['h72A2]=8'h00; mem['h72A3]=8'h00;
    mem['h72A4]=8'h00; mem['h72A5]=8'h00; mem['h72A6]=8'h00; mem['h72A7]=8'h00;
    mem['h72A8]=8'h00; mem['h72A9]=8'h00; mem['h72AA]=8'h00; mem['h72AB]=8'h00;
    mem['h72AC]=8'h00; mem['h72AD]=8'h00; mem['h72AE]=8'h00; mem['h72AF]=8'h00;
    mem['h72B0]=8'h00; mem['h72B1]=8'h00; mem['h72B2]=8'h00; mem['h72B3]=8'h00;
    mem['h72B4]=8'h00; mem['h72B5]=8'h00; mem['h72B6]=8'h00; mem['h72B7]=8'h00;
    mem['h72B8]=8'h00; mem['h72B9]=8'h00; mem['h72BA]=8'h00; mem['h72BB]=8'h00;
    mem['h72BC]=8'h00; mem['h72BD]=8'h00; mem['h72BE]=8'h00; mem['h72BF]=8'h00;
    mem['h72C0]=8'h00; mem['h72C1]=8'h00; mem['h72C2]=8'h00; mem['h72C3]=8'h00;
    mem['h72C4]=8'h00; mem['h72C5]=8'h00; mem['h72C6]=8'h00; mem['h72C7]=8'h00;
    mem['h72C8]=8'h00; mem['h72C9]=8'h00; mem['h72CA]=8'h00; mem['h72CB]=8'h00;
    mem['h72CC]=8'h00; mem['h72CD]=8'h00; mem['h72CE]=8'h00; mem['h72CF]=8'h00;
    mem['h72D0]=8'h00; mem['h72D1]=8'h00; mem['h72D2]=8'h00; mem['h72D3]=8'h00;
    mem['h72D4]=8'h00; mem['h72D5]=8'h00; mem['h72D6]=8'h00; mem['h72D7]=8'h00;
    mem['h72D8]=8'h00; mem['h72D9]=8'h00; mem['h72DA]=8'h00; mem['h72DB]=8'h00;
    mem['h72DC]=8'h00; mem['h72DD]=8'h00; mem['h72DE]=8'h00; mem['h72DF]=8'h00;
    mem['h72E0]=8'h00; mem['h72E1]=8'h00; mem['h72E2]=8'h00; mem['h72E3]=8'h00;
    mem['h72E4]=8'h00; mem['h72E5]=8'h00; mem['h72E6]=8'h00; mem['h72E7]=8'h00;
    mem['h72E8]=8'h00; mem['h72E9]=8'h00; mem['h72EA]=8'h00; mem['h72EB]=8'h00;
    mem['h72EC]=8'h00; mem['h72ED]=8'h00; mem['h72EE]=8'h00; mem['h72EF]=8'h00;
    mem['h72F0]=8'h00; mem['h72F1]=8'h00; mem['h72F2]=8'h00; mem['h72F3]=8'h00;
    mem['h72F4]=8'h00; mem['h72F5]=8'h00; mem['h72F6]=8'h00; mem['h72F7]=8'h00;
    mem['h72F8]=8'h00; mem['h72F9]=8'h00; mem['h72FA]=8'h00; mem['h72FB]=8'h00;
    mem['h72FC]=8'h00; mem['h72FD]=8'h00; mem['h72FE]=8'h00; mem['h72FF]=8'h00;
    mem['h7300]=8'h00; mem['h7301]=8'h00; mem['h7302]=8'h00; mem['h7303]=8'h00;
    mem['h7304]=8'h00; mem['h7305]=8'h00; mem['h7306]=8'h00; mem['h7307]=8'h00;
    mem['h7308]=8'h00; mem['h7309]=8'h00; mem['h730A]=8'h00; mem['h730B]=8'h00;
    mem['h730C]=8'h00; mem['h730D]=8'h00; mem['h730E]=8'h00; mem['h730F]=8'h00;
    mem['h7310]=8'h00; mem['h7311]=8'h00; mem['h7312]=8'h00; mem['h7313]=8'h00;
    mem['h7314]=8'h00; mem['h7315]=8'h00; mem['h7316]=8'h00; mem['h7317]=8'h00;
    mem['h7318]=8'h00; mem['h7319]=8'h00; mem['h731A]=8'h00; mem['h731B]=8'h00;
    mem['h731C]=8'h00; mem['h731D]=8'h00; mem['h731E]=8'h00; mem['h731F]=8'h00;
    mem['h7320]=8'h00; mem['h7321]=8'h00; mem['h7322]=8'h00; mem['h7323]=8'h00;
    mem['h7324]=8'h00; mem['h7325]=8'h00; mem['h7326]=8'h00; mem['h7327]=8'h00;
    mem['h7328]=8'h00; mem['h7329]=8'h00; mem['h732A]=8'h00; mem['h732B]=8'h00;
    mem['h732C]=8'h00; mem['h732D]=8'h00; mem['h732E]=8'h00; mem['h732F]=8'h00;
    mem['h7330]=8'h00; mem['h7331]=8'h00; mem['h7332]=8'h00; mem['h7333]=8'h00;
    mem['h7334]=8'h00; mem['h7335]=8'h00; mem['h7336]=8'h00; mem['h7337]=8'h00;
    mem['h7338]=8'h00; mem['h7339]=8'h00; mem['h733A]=8'h00; mem['h733B]=8'h00;
    mem['h733C]=8'h00; mem['h733D]=8'h00; mem['h733E]=8'h00; mem['h733F]=8'h00;
    mem['h7340]=8'h00; mem['h7341]=8'h00; mem['h7342]=8'h00; mem['h7343]=8'h00;
    mem['h7344]=8'h00; mem['h7345]=8'h00; mem['h7346]=8'h00; mem['h7347]=8'h00;
    mem['h7348]=8'h00; mem['h7349]=8'h00; mem['h734A]=8'h00; mem['h734B]=8'h00;
    mem['h734C]=8'h00; mem['h734D]=8'h00; mem['h734E]=8'h00; mem['h734F]=8'h00;
    mem['h7350]=8'h00; mem['h7351]=8'h00; mem['h7352]=8'h00; mem['h7353]=8'h00;
    mem['h7354]=8'h00; mem['h7355]=8'h00; mem['h7356]=8'h00; mem['h7357]=8'h00;
    mem['h7358]=8'h00; mem['h7359]=8'h00; mem['h735A]=8'h00; mem['h735B]=8'h00;
    mem['h735C]=8'h00; mem['h735D]=8'h00; mem['h735E]=8'h00; mem['h735F]=8'h00;
    mem['h7360]=8'h00; mem['h7361]=8'h00; mem['h7362]=8'h00; mem['h7363]=8'h00;
    mem['h7364]=8'h00; mem['h7365]=8'h00; mem['h7366]=8'h00; mem['h7367]=8'h00;
    mem['h7368]=8'h00; mem['h7369]=8'h00; mem['h736A]=8'h00; mem['h736B]=8'h00;
    mem['h736C]=8'h00; mem['h736D]=8'h00; mem['h736E]=8'h00; mem['h736F]=8'h00;
    mem['h7370]=8'h00; mem['h7371]=8'h00; mem['h7372]=8'h00; mem['h7373]=8'h00;
    mem['h7374]=8'h00; mem['h7375]=8'h00; mem['h7376]=8'h00; mem['h7377]=8'h00;
    mem['h7378]=8'h00; mem['h7379]=8'h00; mem['h737A]=8'h00; mem['h737B]=8'h00;
    mem['h737C]=8'h00; mem['h737D]=8'h00; mem['h737E]=8'h00; mem['h737F]=8'h00;
    mem['h7380]=8'h00; mem['h7381]=8'h00; mem['h7382]=8'h00; mem['h7383]=8'h00;
    mem['h7384]=8'h00; mem['h7385]=8'h00; mem['h7386]=8'h00; mem['h7387]=8'h00;
    mem['h7388]=8'h00; mem['h7389]=8'h00; mem['h738A]=8'h00; mem['h738B]=8'h00;
    mem['h738C]=8'h00; mem['h738D]=8'h00; mem['h738E]=8'h00; mem['h738F]=8'h00;
    mem['h7390]=8'h00; mem['h7391]=8'h00; mem['h7392]=8'h00; mem['h7393]=8'h00;
    mem['h7394]=8'h00; mem['h7395]=8'h00; mem['h7396]=8'h00; mem['h7397]=8'h00;
    mem['h7398]=8'h00; mem['h7399]=8'h00; mem['h739A]=8'h00; mem['h739B]=8'h00;
    mem['h739C]=8'h00; mem['h739D]=8'h00; mem['h739E]=8'h00; mem['h739F]=8'h00;
    mem['h73A0]=8'h00; mem['h73A1]=8'h00; mem['h73A2]=8'h00; mem['h73A3]=8'h00;
    mem['h73A4]=8'h00; mem['h73A5]=8'h00; mem['h73A6]=8'h00; mem['h73A7]=8'h00;
    mem['h73A8]=8'h00; mem['h73A9]=8'h00; mem['h73AA]=8'h00; mem['h73AB]=8'h00;
    mem['h73AC]=8'h00; mem['h73AD]=8'h00; mem['h73AE]=8'h00; mem['h73AF]=8'h00;
    mem['h73B0]=8'h00; mem['h73B1]=8'h00; mem['h73B2]=8'h00; mem['h73B3]=8'h00;
    mem['h73B4]=8'h00; mem['h73B5]=8'h00; mem['h73B6]=8'h00; mem['h73B7]=8'h00;
    mem['h73B8]=8'h00; mem['h73B9]=8'h00; mem['h73BA]=8'h00; mem['h73BB]=8'h00;
    mem['h73BC]=8'h00; mem['h73BD]=8'h00; mem['h73BE]=8'h00; mem['h73BF]=8'h00;
    mem['h73C0]=8'h00; mem['h73C1]=8'h00; mem['h73C2]=8'h00; mem['h73C3]=8'h00;
    mem['h73C4]=8'h00; mem['h73C5]=8'h00; mem['h73C6]=8'h00; mem['h73C7]=8'h00;
    mem['h73C8]=8'h00; mem['h73C9]=8'h00; mem['h73CA]=8'h00; mem['h73CB]=8'h00;
    mem['h73CC]=8'h00; mem['h73CD]=8'h00; mem['h73CE]=8'h00; mem['h73CF]=8'h00;
    mem['h73D0]=8'h00; mem['h73D1]=8'h00; mem['h73D2]=8'h00; mem['h73D3]=8'h00;
    mem['h73D4]=8'h00; mem['h73D5]=8'h00; mem['h73D6]=8'h00; mem['h73D7]=8'h00;
    mem['h73D8]=8'h00; mem['h73D9]=8'h00; mem['h73DA]=8'h00; mem['h73DB]=8'h00;
    mem['h73DC]=8'h00; mem['h73DD]=8'h00; mem['h73DE]=8'h00; mem['h73DF]=8'h00;
    mem['h73E0]=8'h00; mem['h73E1]=8'h00; mem['h73E2]=8'h00; mem['h73E3]=8'h00;
    mem['h73E4]=8'h00; mem['h73E5]=8'h00; mem['h73E6]=8'h00; mem['h73E7]=8'h00;
    mem['h73E8]=8'h00; mem['h73E9]=8'h00; mem['h73EA]=8'h00; mem['h73EB]=8'h00;
    mem['h73EC]=8'h00; mem['h73ED]=8'h00; mem['h73EE]=8'h00; mem['h73EF]=8'h00;
    mem['h73F0]=8'h00; mem['h73F1]=8'h00; mem['h73F2]=8'h00; mem['h73F3]=8'h00;
    mem['h73F4]=8'h00; mem['h73F5]=8'h00; mem['h73F6]=8'h00; mem['h73F7]=8'h00;
    mem['h73F8]=8'h00; mem['h73F9]=8'h00; mem['h73FA]=8'h00; mem['h73FB]=8'h00;
    mem['h73FC]=8'h00; mem['h73FD]=8'h00; mem['h73FE]=8'h00; mem['h73FF]=8'h00;
    mem['h7400]=8'h00; mem['h7401]=8'h00; mem['h7402]=8'h00; mem['h7403]=8'h00;
    mem['h7404]=8'h00; mem['h7405]=8'h00; mem['h7406]=8'h00; mem['h7407]=8'h00;
    mem['h7408]=8'h00; mem['h7409]=8'h00; mem['h740A]=8'h00; mem['h740B]=8'h00;
    mem['h740C]=8'h00; mem['h740D]=8'h00; mem['h740E]=8'h00; mem['h740F]=8'h00;
    mem['h7410]=8'h00; mem['h7411]=8'h00; mem['h7412]=8'h00; mem['h7413]=8'h00;
    mem['h7414]=8'h00; mem['h7415]=8'h00; mem['h7416]=8'h00; mem['h7417]=8'h00;
    mem['h7418]=8'h00; mem['h7419]=8'h00; mem['h741A]=8'h00; mem['h741B]=8'h00;
    mem['h741C]=8'h00; mem['h741D]=8'h00; mem['h741E]=8'h00; mem['h741F]=8'h00;
    mem['h7420]=8'h00; mem['h7421]=8'h00; mem['h7422]=8'h00; mem['h7423]=8'h00;
    mem['h7424]=8'h00; mem['h7425]=8'h00; mem['h7426]=8'h00; mem['h7427]=8'h00;
    mem['h7428]=8'h00; mem['h7429]=8'h00; mem['h742A]=8'h00; mem['h742B]=8'h00;
    mem['h742C]=8'h00; mem['h742D]=8'h00; mem['h742E]=8'h00; mem['h742F]=8'h00;
    mem['h7430]=8'h00; mem['h7431]=8'h00; mem['h7432]=8'h00; mem['h7433]=8'h00;
    mem['h7434]=8'h00; mem['h7435]=8'h00; mem['h7436]=8'h00; mem['h7437]=8'h00;
    mem['h7438]=8'h00; mem['h7439]=8'h00; mem['h743A]=8'h00; mem['h743B]=8'h00;
    mem['h743C]=8'h00; mem['h743D]=8'h00; mem['h743E]=8'h00; mem['h743F]=8'h00;
    mem['h7440]=8'h00; mem['h7441]=8'h00; mem['h7442]=8'h00; mem['h7443]=8'h00;
    mem['h7444]=8'h00; mem['h7445]=8'h00; mem['h7446]=8'h00; mem['h7447]=8'h00;
    mem['h7448]=8'h00; mem['h7449]=8'h00; mem['h744A]=8'h00; mem['h744B]=8'h00;
    mem['h744C]=8'h00; mem['h744D]=8'h00; mem['h744E]=8'h00; mem['h744F]=8'h00;
    mem['h7450]=8'h00; mem['h7451]=8'h00; mem['h7452]=8'h00; mem['h7453]=8'h00;
    mem['h7454]=8'h00; mem['h7455]=8'h00; mem['h7456]=8'h00; mem['h7457]=8'h00;
    mem['h7458]=8'h00; mem['h7459]=8'h00; mem['h745A]=8'h00; mem['h745B]=8'h00;
    mem['h745C]=8'h00; mem['h745D]=8'h00; mem['h745E]=8'h00; mem['h745F]=8'h00;
    mem['h7460]=8'h00; mem['h7461]=8'h00; mem['h7462]=8'h00; mem['h7463]=8'h00;
    mem['h7464]=8'h00; mem['h7465]=8'h00; mem['h7466]=8'h00; mem['h7467]=8'h00;
    mem['h7468]=8'h00; mem['h7469]=8'h00; mem['h746A]=8'h00; mem['h746B]=8'h00;
    mem['h746C]=8'h00; mem['h746D]=8'h00; mem['h746E]=8'h00; mem['h746F]=8'h00;
    mem['h7470]=8'h00; mem['h7471]=8'h00; mem['h7472]=8'h00; mem['h7473]=8'h00;
    mem['h7474]=8'h00; mem['h7475]=8'h00; mem['h7476]=8'h00; mem['h7477]=8'h00;
    mem['h7478]=8'h00; mem['h7479]=8'h00; mem['h747A]=8'h00; mem['h747B]=8'h00;
    mem['h747C]=8'h00; mem['h747D]=8'h00; mem['h747E]=8'h00; mem['h747F]=8'h00;
    mem['h7480]=8'h00; mem['h7481]=8'h00; mem['h7482]=8'h00; mem['h7483]=8'h00;
    mem['h7484]=8'h00; mem['h7485]=8'h00; mem['h7486]=8'h00; mem['h7487]=8'h00;
    mem['h7488]=8'h00; mem['h7489]=8'h00; mem['h748A]=8'h00; mem['h748B]=8'h00;
    mem['h748C]=8'h00; mem['h748D]=8'h00; mem['h748E]=8'h00; mem['h748F]=8'h00;
    mem['h7490]=8'h00; mem['h7491]=8'h00; mem['h7492]=8'h00; mem['h7493]=8'h00;
    mem['h7494]=8'h00; mem['h7495]=8'h00; mem['h7496]=8'h00; mem['h7497]=8'h00;
    mem['h7498]=8'h00; mem['h7499]=8'h00; mem['h749A]=8'h00; mem['h749B]=8'h00;
    mem['h749C]=8'h00; mem['h749D]=8'h00; mem['h749E]=8'h00; mem['h749F]=8'h00;
    mem['h74A0]=8'h00; mem['h74A1]=8'h00; mem['h74A2]=8'h00; mem['h74A3]=8'h00;
    mem['h74A4]=8'h00; mem['h74A5]=8'h00; mem['h74A6]=8'h00; mem['h74A7]=8'h00;
    mem['h74A8]=8'h00; mem['h74A9]=8'h00; mem['h74AA]=8'h00; mem['h74AB]=8'h00;
    mem['h74AC]=8'h00; mem['h74AD]=8'h00; mem['h74AE]=8'h00; mem['h74AF]=8'h00;
    mem['h74B0]=8'h00; mem['h74B1]=8'h00; mem['h74B2]=8'h00; mem['h74B3]=8'h00;
    mem['h74B4]=8'h00; mem['h74B5]=8'h00; mem['h74B6]=8'h00; mem['h74B7]=8'h00;
    mem['h74B8]=8'h00; mem['h74B9]=8'h00; mem['h74BA]=8'h00; mem['h74BB]=8'h00;
    mem['h74BC]=8'h00; mem['h74BD]=8'h00; mem['h74BE]=8'h00; mem['h74BF]=8'h00;
    mem['h74C0]=8'h00; mem['h74C1]=8'h00; mem['h74C2]=8'h00; mem['h74C3]=8'h00;
    mem['h74C4]=8'h00; mem['h74C5]=8'h00; mem['h74C6]=8'h00; mem['h74C7]=8'h00;
    mem['h74C8]=8'h00; mem['h74C9]=8'h00; mem['h74CA]=8'h00; mem['h74CB]=8'h00;
    mem['h74CC]=8'h00; mem['h74CD]=8'h00; mem['h74CE]=8'h00; mem['h74CF]=8'h00;
    mem['h74D0]=8'h00; mem['h74D1]=8'h00; mem['h74D2]=8'h00; mem['h74D3]=8'h00;
    mem['h74D4]=8'h00; mem['h74D5]=8'h00; mem['h74D6]=8'h00; mem['h74D7]=8'h00;
    mem['h74D8]=8'h00; mem['h74D9]=8'h00; mem['h74DA]=8'h00; mem['h74DB]=8'h00;
    mem['h74DC]=8'h00; mem['h74DD]=8'h00; mem['h74DE]=8'h00; mem['h74DF]=8'h00;
    mem['h74E0]=8'h00; mem['h74E1]=8'h00; mem['h74E2]=8'h00; mem['h74E3]=8'h00;
    mem['h74E4]=8'h00; mem['h74E5]=8'h00; mem['h74E6]=8'h00; mem['h74E7]=8'h00;
    mem['h74E8]=8'h00; mem['h74E9]=8'h00; mem['h74EA]=8'h00; mem['h74EB]=8'h00;
    mem['h74EC]=8'h00; mem['h74ED]=8'h00; mem['h74EE]=8'h00; mem['h74EF]=8'h00;
    mem['h74F0]=8'h00; mem['h74F1]=8'h00; mem['h74F2]=8'h00; mem['h74F3]=8'h00;
    mem['h74F4]=8'h00; mem['h74F5]=8'h00; mem['h74F6]=8'h00; mem['h74F7]=8'h00;
    mem['h74F8]=8'h00; mem['h74F9]=8'h00; mem['h74FA]=8'h00; mem['h74FB]=8'h00;
    mem['h74FC]=8'h00; mem['h74FD]=8'h00; mem['h74FE]=8'h00; mem['h74FF]=8'h00;
    mem['h7500]=8'h00; mem['h7501]=8'h00; mem['h7502]=8'h00; mem['h7503]=8'h00;
    mem['h7504]=8'h00; mem['h7505]=8'h00; mem['h7506]=8'h00; mem['h7507]=8'h00;
    mem['h7508]=8'h00; mem['h7509]=8'h00; mem['h750A]=8'h00; mem['h750B]=8'h00;
    mem['h750C]=8'h00; mem['h750D]=8'h00; mem['h750E]=8'h00; mem['h750F]=8'h00;
    mem['h7510]=8'h00; mem['h7511]=8'h00; mem['h7512]=8'h00; mem['h7513]=8'h00;
    mem['h7514]=8'h00; mem['h7515]=8'h00; mem['h7516]=8'h00; mem['h7517]=8'h00;
    mem['h7518]=8'h00; mem['h7519]=8'h00; mem['h751A]=8'h00; mem['h751B]=8'h00;
    mem['h751C]=8'h00; mem['h751D]=8'h00; mem['h751E]=8'h00; mem['h751F]=8'h00;
    mem['h7520]=8'h00; mem['h7521]=8'h00; mem['h7522]=8'h00; mem['h7523]=8'h00;
    mem['h7524]=8'h00; mem['h7525]=8'h00; mem['h7526]=8'h00; mem['h7527]=8'h00;
    mem['h7528]=8'h00; mem['h7529]=8'h00; mem['h752A]=8'h00; mem['h752B]=8'h00;
    mem['h752C]=8'h00; mem['h752D]=8'h00; mem['h752E]=8'h00; mem['h752F]=8'h00;
    mem['h7530]=8'h00; mem['h7531]=8'h00; mem['h7532]=8'h00; mem['h7533]=8'h00;
    mem['h7534]=8'h00; mem['h7535]=8'h00; mem['h7536]=8'h00; mem['h7537]=8'h00;
    mem['h7538]=8'h00; mem['h7539]=8'h00; mem['h753A]=8'h00; mem['h753B]=8'h00;
    mem['h753C]=8'h00; mem['h753D]=8'h00; mem['h753E]=8'h00; mem['h753F]=8'h00;
    mem['h7540]=8'h00; mem['h7541]=8'h00; mem['h7542]=8'h00; mem['h7543]=8'h00;
    mem['h7544]=8'h00; mem['h7545]=8'h00; mem['h7546]=8'h00; mem['h7547]=8'h00;
    mem['h7548]=8'h00; mem['h7549]=8'h00; mem['h754A]=8'h00; mem['h754B]=8'h00;
    mem['h754C]=8'h00; mem['h754D]=8'h00; mem['h754E]=8'h00; mem['h754F]=8'h00;
    mem['h7550]=8'h00; mem['h7551]=8'h00; mem['h7552]=8'h00; mem['h7553]=8'h00;
    mem['h7554]=8'h00; mem['h7555]=8'h00; mem['h7556]=8'h00; mem['h7557]=8'h00;
    mem['h7558]=8'h00; mem['h7559]=8'h00; mem['h755A]=8'h00; mem['h755B]=8'h00;
    mem['h755C]=8'h00; mem['h755D]=8'h00; mem['h755E]=8'h00; mem['h755F]=8'h00;
    mem['h7560]=8'h00; mem['h7561]=8'h00; mem['h7562]=8'h00; mem['h7563]=8'h00;
    mem['h7564]=8'h00; mem['h7565]=8'h00; mem['h7566]=8'h00; mem['h7567]=8'h00;
    mem['h7568]=8'h00; mem['h7569]=8'h00; mem['h756A]=8'h00; mem['h756B]=8'h00;
    mem['h756C]=8'h00; mem['h756D]=8'h00; mem['h756E]=8'h00; mem['h756F]=8'h00;
    mem['h7570]=8'h00; mem['h7571]=8'h00; mem['h7572]=8'h00; mem['h7573]=8'h00;
    mem['h7574]=8'h00; mem['h7575]=8'h00; mem['h7576]=8'h00; mem['h7577]=8'h00;
    mem['h7578]=8'h00; mem['h7579]=8'h00; mem['h757A]=8'h00; mem['h757B]=8'h00;
    mem['h757C]=8'h00; mem['h757D]=8'h00; mem['h757E]=8'h00; mem['h757F]=8'h00;
    mem['h7580]=8'h00; mem['h7581]=8'h00; mem['h7582]=8'h00; mem['h7583]=8'h00;
    mem['h7584]=8'h00; mem['h7585]=8'h00; mem['h7586]=8'h00; mem['h7587]=8'h00;
    mem['h7588]=8'h00; mem['h7589]=8'h00; mem['h758A]=8'h00; mem['h758B]=8'h00;
    mem['h758C]=8'h00; mem['h758D]=8'h00; mem['h758E]=8'h00; mem['h758F]=8'h00;
    mem['h7590]=8'h00; mem['h7591]=8'h00; mem['h7592]=8'h00; mem['h7593]=8'h00;
    mem['h7594]=8'h00; mem['h7595]=8'h00; mem['h7596]=8'h00; mem['h7597]=8'h00;
    mem['h7598]=8'h00; mem['h7599]=8'h00; mem['h759A]=8'h00; mem['h759B]=8'h00;
    mem['h759C]=8'h00; mem['h759D]=8'h00; mem['h759E]=8'h00; mem['h759F]=8'h00;
    mem['h75A0]=8'h00; mem['h75A1]=8'h00; mem['h75A2]=8'h00; mem['h75A3]=8'h00;
    mem['h75A4]=8'h00; mem['h75A5]=8'h00; mem['h75A6]=8'h00; mem['h75A7]=8'h00;
    mem['h75A8]=8'h00; mem['h75A9]=8'h00; mem['h75AA]=8'h00; mem['h75AB]=8'h00;
    mem['h75AC]=8'h00; mem['h75AD]=8'h00; mem['h75AE]=8'h00; mem['h75AF]=8'h00;
    mem['h75B0]=8'h00; mem['h75B1]=8'h00; mem['h75B2]=8'h00; mem['h75B3]=8'h00;
    mem['h75B4]=8'h00; mem['h75B5]=8'h00; mem['h75B6]=8'h00; mem['h75B7]=8'h00;
    mem['h75B8]=8'h00; mem['h75B9]=8'h00; mem['h75BA]=8'h00; mem['h75BB]=8'h00;
    mem['h75BC]=8'h00; mem['h75BD]=8'h00; mem['h75BE]=8'h00; mem['h75BF]=8'h00;
    mem['h75C0]=8'h00; mem['h75C1]=8'h00; mem['h75C2]=8'h00; mem['h75C3]=8'h00;
    mem['h75C4]=8'h00; mem['h75C5]=8'h00; mem['h75C6]=8'h00; mem['h75C7]=8'h00;
    mem['h75C8]=8'h00; mem['h75C9]=8'h00; mem['h75CA]=8'h00; mem['h75CB]=8'h00;
    mem['h75CC]=8'h00; mem['h75CD]=8'h00; mem['h75CE]=8'h00; mem['h75CF]=8'h00;
    mem['h75D0]=8'h00; mem['h75D1]=8'h00; mem['h75D2]=8'h00; mem['h75D3]=8'h00;
    mem['h75D4]=8'h00; mem['h75D5]=8'h00; mem['h75D6]=8'h00; mem['h75D7]=8'h00;
    mem['h75D8]=8'h00; mem['h75D9]=8'h00; mem['h75DA]=8'h00; mem['h75DB]=8'h00;
    mem['h75DC]=8'h00; mem['h75DD]=8'h00; mem['h75DE]=8'h00; mem['h75DF]=8'h00;
    mem['h75E0]=8'h00; mem['h75E1]=8'h00; mem['h75E2]=8'h00; mem['h75E3]=8'h00;
    mem['h75E4]=8'h00; mem['h75E5]=8'h00; mem['h75E6]=8'h00; mem['h75E7]=8'h00;
    mem['h75E8]=8'h00; mem['h75E9]=8'h00; mem['h75EA]=8'h00; mem['h75EB]=8'h00;
    mem['h75EC]=8'h00; mem['h75ED]=8'h00; mem['h75EE]=8'h00; mem['h75EF]=8'h00;
    mem['h75F0]=8'h00; mem['h75F1]=8'h00; mem['h75F2]=8'h00; mem['h75F3]=8'h00;
    mem['h75F4]=8'h00; mem['h75F5]=8'h00; mem['h75F6]=8'h00; mem['h75F7]=8'h00;
    mem['h75F8]=8'h00; mem['h75F9]=8'h00; mem['h75FA]=8'h00; mem['h75FB]=8'h00;
    mem['h75FC]=8'h00; mem['h75FD]=8'h00; mem['h75FE]=8'h00; mem['h75FF]=8'h00;
    mem['h7600]=8'h00; mem['h7601]=8'h00; mem['h7602]=8'h00; mem['h7603]=8'h00;
    mem['h7604]=8'h00; mem['h7605]=8'h00; mem['h7606]=8'h00; mem['h7607]=8'h00;
    mem['h7608]=8'h00; mem['h7609]=8'h00; mem['h760A]=8'h00; mem['h760B]=8'h00;
    mem['h760C]=8'h00; mem['h760D]=8'h00; mem['h760E]=8'h00; mem['h760F]=8'h00;
    mem['h7610]=8'h00; mem['h7611]=8'h00; mem['h7612]=8'h00; mem['h7613]=8'h00;
    mem['h7614]=8'h00; mem['h7615]=8'h00; mem['h7616]=8'h00; mem['h7617]=8'h00;
    mem['h7618]=8'h00; mem['h7619]=8'h00; mem['h761A]=8'h00; mem['h761B]=8'h00;
    mem['h761C]=8'h00; mem['h761D]=8'h00; mem['h761E]=8'h00; mem['h761F]=8'h00;
    mem['h7620]=8'h00; mem['h7621]=8'h00; mem['h7622]=8'h00; mem['h7623]=8'h00;
    mem['h7624]=8'h00; mem['h7625]=8'h00; mem['h7626]=8'h00; mem['h7627]=8'h00;
    mem['h7628]=8'h00; mem['h7629]=8'h00; mem['h762A]=8'h00; mem['h762B]=8'h00;
    mem['h762C]=8'h00; mem['h762D]=8'h00; mem['h762E]=8'h00; mem['h762F]=8'h00;
    mem['h7630]=8'h00; mem['h7631]=8'h00; mem['h7632]=8'h00; mem['h7633]=8'h00;
    mem['h7634]=8'h00; mem['h7635]=8'h00; mem['h7636]=8'h00; mem['h7637]=8'h00;
    mem['h7638]=8'h00; mem['h7639]=8'h00; mem['h763A]=8'h00; mem['h763B]=8'h00;
    mem['h763C]=8'h00; mem['h763D]=8'h00; mem['h763E]=8'h00; mem['h763F]=8'h00;
    mem['h7640]=8'h00; mem['h7641]=8'h00; mem['h7642]=8'h00; mem['h7643]=8'h00;
    mem['h7644]=8'h00; mem['h7645]=8'h00; mem['h7646]=8'h00; mem['h7647]=8'h00;
    mem['h7648]=8'h00; mem['h7649]=8'h00; mem['h764A]=8'h00; mem['h764B]=8'h00;
    mem['h764C]=8'h00; mem['h764D]=8'h00; mem['h764E]=8'h00; mem['h764F]=8'h00;
    mem['h7650]=8'h00; mem['h7651]=8'h00; mem['h7652]=8'h00; mem['h7653]=8'h00;
    mem['h7654]=8'h00; mem['h7655]=8'h00; mem['h7656]=8'h00; mem['h7657]=8'h00;
    mem['h7658]=8'h00; mem['h7659]=8'h00; mem['h765A]=8'h00; mem['h765B]=8'h00;
    mem['h765C]=8'h00; mem['h765D]=8'h00; mem['h765E]=8'h00; mem['h765F]=8'h00;
    mem['h7660]=8'h00; mem['h7661]=8'h00; mem['h7662]=8'h00; mem['h7663]=8'h00;
    mem['h7664]=8'h00; mem['h7665]=8'h00; mem['h7666]=8'h00; mem['h7667]=8'h00;
    mem['h7668]=8'h00; mem['h7669]=8'h00; mem['h766A]=8'h00; mem['h766B]=8'h00;
    mem['h766C]=8'h00; mem['h766D]=8'h00; mem['h766E]=8'h00; mem['h766F]=8'h00;
    mem['h7670]=8'h00; mem['h7671]=8'h00; mem['h7672]=8'h00; mem['h7673]=8'h00;
    mem['h7674]=8'h00; mem['h7675]=8'h00; mem['h7676]=8'h00; mem['h7677]=8'h00;
    mem['h7678]=8'h00; mem['h7679]=8'h00; mem['h767A]=8'h00; mem['h767B]=8'h00;
    mem['h767C]=8'h00; mem['h767D]=8'h00; mem['h767E]=8'h00; mem['h767F]=8'h00;
    mem['h7680]=8'h00; mem['h7681]=8'h00; mem['h7682]=8'h00; mem['h7683]=8'h00;
    mem['h7684]=8'h00; mem['h7685]=8'h00; mem['h7686]=8'h00; mem['h7687]=8'h00;
    mem['h7688]=8'h00; mem['h7689]=8'h00; mem['h768A]=8'h00; mem['h768B]=8'h00;
    mem['h768C]=8'h00; mem['h768D]=8'h00; mem['h768E]=8'h00; mem['h768F]=8'h00;
    mem['h7690]=8'h00; mem['h7691]=8'h00; mem['h7692]=8'h00; mem['h7693]=8'h00;
    mem['h7694]=8'h00; mem['h7695]=8'h00; mem['h7696]=8'h00; mem['h7697]=8'h00;
    mem['h7698]=8'h00; mem['h7699]=8'h00; mem['h769A]=8'h00; mem['h769B]=8'h00;
    mem['h769C]=8'h00; mem['h769D]=8'h00; mem['h769E]=8'h00; mem['h769F]=8'h00;
    mem['h76A0]=8'h00; mem['h76A1]=8'h00; mem['h76A2]=8'h00; mem['h76A3]=8'h00;
    mem['h76A4]=8'h00; mem['h76A5]=8'h00; mem['h76A6]=8'h00; mem['h76A7]=8'h00;
    mem['h76A8]=8'h00; mem['h76A9]=8'h00; mem['h76AA]=8'h00; mem['h76AB]=8'h00;
    mem['h76AC]=8'h00; mem['h76AD]=8'h00; mem['h76AE]=8'h00; mem['h76AF]=8'h00;
    mem['h76B0]=8'h00; mem['h76B1]=8'h00; mem['h76B2]=8'h00; mem['h76B3]=8'h00;
    mem['h76B4]=8'h00; mem['h76B5]=8'h00; mem['h76B6]=8'h00; mem['h76B7]=8'h00;
    mem['h76B8]=8'h00; mem['h76B9]=8'h00; mem['h76BA]=8'h00; mem['h76BB]=8'h00;
    mem['h76BC]=8'h00; mem['h76BD]=8'h00; mem['h76BE]=8'h00; mem['h76BF]=8'h00;
    mem['h76C0]=8'h00; mem['h76C1]=8'h00; mem['h76C2]=8'h00; mem['h76C3]=8'h00;
    mem['h76C4]=8'h00; mem['h76C5]=8'h00; mem['h76C6]=8'h00; mem['h76C7]=8'h00;
    mem['h76C8]=8'h00; mem['h76C9]=8'h00; mem['h76CA]=8'h00; mem['h76CB]=8'h00;
    mem['h76CC]=8'h00; mem['h76CD]=8'h00; mem['h76CE]=8'h00; mem['h76CF]=8'h00;
    mem['h76D0]=8'h00; mem['h76D1]=8'h00; mem['h76D2]=8'h00; mem['h76D3]=8'h00;
    mem['h76D4]=8'h00; mem['h76D5]=8'h00; mem['h76D6]=8'h00; mem['h76D7]=8'h00;
    mem['h76D8]=8'h00; mem['h76D9]=8'h00; mem['h76DA]=8'h00; mem['h76DB]=8'h00;
    mem['h76DC]=8'h00; mem['h76DD]=8'h00; mem['h76DE]=8'h00; mem['h76DF]=8'h00;
    mem['h76E0]=8'h00; mem['h76E1]=8'h00; mem['h76E2]=8'h00; mem['h76E3]=8'h00;
    mem['h76E4]=8'h00; mem['h76E5]=8'h00; mem['h76E6]=8'h00; mem['h76E7]=8'h00;
    mem['h76E8]=8'h00; mem['h76E9]=8'h00; mem['h76EA]=8'h00; mem['h76EB]=8'h00;
    mem['h76EC]=8'h00; mem['h76ED]=8'h00; mem['h76EE]=8'h00; mem['h76EF]=8'h00;
    mem['h76F0]=8'h00; mem['h76F1]=8'h00; mem['h76F2]=8'h00; mem['h76F3]=8'h00;
    mem['h76F4]=8'h00; mem['h76F5]=8'h00; mem['h76F6]=8'h00; mem['h76F7]=8'h00;
    mem['h76F8]=8'h00; mem['h76F9]=8'h00; mem['h76FA]=8'h00; mem['h76FB]=8'h00;
    mem['h76FC]=8'h00; mem['h76FD]=8'h00; mem['h76FE]=8'h00; mem['h76FF]=8'h00;
    mem['h7700]=8'h00; mem['h7701]=8'h00; mem['h7702]=8'h00; mem['h7703]=8'h00;
    mem['h7704]=8'h00; mem['h7705]=8'h00; mem['h7706]=8'h00; mem['h7707]=8'h00;
    mem['h7708]=8'h00; mem['h7709]=8'h00; mem['h770A]=8'h00; mem['h770B]=8'h00;
    mem['h770C]=8'h00; mem['h770D]=8'h00; mem['h770E]=8'h00; mem['h770F]=8'h00;
    mem['h7710]=8'h00; mem['h7711]=8'h00; mem['h7712]=8'h00; mem['h7713]=8'h00;
    mem['h7714]=8'h00; mem['h7715]=8'h00; mem['h7716]=8'h00; mem['h7717]=8'h00;
    mem['h7718]=8'h00; mem['h7719]=8'h00; mem['h771A]=8'h00; mem['h771B]=8'h00;
    mem['h771C]=8'h00; mem['h771D]=8'h00; mem['h771E]=8'h00; mem['h771F]=8'h00;
    mem['h7720]=8'h00; mem['h7721]=8'h00; mem['h7722]=8'h00; mem['h7723]=8'h00;
    mem['h7724]=8'h00; mem['h7725]=8'h00; mem['h7726]=8'h00; mem['h7727]=8'h00;
    mem['h7728]=8'h00; mem['h7729]=8'h00; mem['h772A]=8'h00; mem['h772B]=8'h00;
    mem['h772C]=8'h00; mem['h772D]=8'h00; mem['h772E]=8'h00; mem['h772F]=8'h00;
    mem['h7730]=8'h00; mem['h7731]=8'h00; mem['h7732]=8'h00; mem['h7733]=8'h00;
    mem['h7734]=8'h00; mem['h7735]=8'h00; mem['h7736]=8'h00; mem['h7737]=8'h00;
    mem['h7738]=8'h00; mem['h7739]=8'h00; mem['h773A]=8'h00; mem['h773B]=8'h00;
    mem['h773C]=8'h00; mem['h773D]=8'h00; mem['h773E]=8'h00; mem['h773F]=8'h00;
    mem['h7740]=8'h00; mem['h7741]=8'h00; mem['h7742]=8'h00; mem['h7743]=8'h00;
    mem['h7744]=8'h00; mem['h7745]=8'h00; mem['h7746]=8'h00; mem['h7747]=8'h00;
    mem['h7748]=8'h00; mem['h7749]=8'h00; mem['h774A]=8'h00; mem['h774B]=8'h00;
    mem['h774C]=8'h00; mem['h774D]=8'h00; mem['h774E]=8'h00; mem['h774F]=8'h00;
    mem['h7750]=8'h00; mem['h7751]=8'h00; mem['h7752]=8'h00; mem['h7753]=8'h00;
    mem['h7754]=8'h00; mem['h7755]=8'h00; mem['h7756]=8'h00; mem['h7757]=8'h00;
    mem['h7758]=8'h00; mem['h7759]=8'h00; mem['h775A]=8'h00; mem['h775B]=8'h00;
    mem['h775C]=8'h00; mem['h775D]=8'h00; mem['h775E]=8'h00; mem['h775F]=8'h00;
    mem['h7760]=8'h00; mem['h7761]=8'h00; mem['h7762]=8'h00; mem['h7763]=8'h00;
    mem['h7764]=8'h00; mem['h7765]=8'h00; mem['h7766]=8'h00; mem['h7767]=8'h00;
    mem['h7768]=8'h00; mem['h7769]=8'h00; mem['h776A]=8'h00; mem['h776B]=8'h00;
    mem['h776C]=8'h00; mem['h776D]=8'h00; mem['h776E]=8'h00; mem['h776F]=8'h00;
    mem['h7770]=8'h00; mem['h7771]=8'h00; mem['h7772]=8'h00; mem['h7773]=8'h00;
    mem['h7774]=8'h00; mem['h7775]=8'h00; mem['h7776]=8'h00; mem['h7777]=8'h00;
    mem['h7778]=8'h00; mem['h7779]=8'h00; mem['h777A]=8'h00; mem['h777B]=8'h00;
    mem['h777C]=8'h00; mem['h777D]=8'h00; mem['h777E]=8'h00; mem['h777F]=8'h00;
    mem['h7780]=8'h00; mem['h7781]=8'h00; mem['h7782]=8'h00; mem['h7783]=8'h00;
    mem['h7784]=8'h00; mem['h7785]=8'h00; mem['h7786]=8'h00; mem['h7787]=8'h00;
    mem['h7788]=8'h00; mem['h7789]=8'h00; mem['h778A]=8'h00; mem['h778B]=8'h00;
    mem['h778C]=8'h00; mem['h778D]=8'h00; mem['h778E]=8'h00; mem['h778F]=8'h00;
    mem['h7790]=8'h00; mem['h7791]=8'h00; mem['h7792]=8'h00; mem['h7793]=8'h00;
    mem['h7794]=8'h00; mem['h7795]=8'h00; mem['h7796]=8'h00; mem['h7797]=8'h00;
    mem['h7798]=8'h00; mem['h7799]=8'h00; mem['h779A]=8'h00; mem['h779B]=8'h00;
    mem['h779C]=8'h00; mem['h779D]=8'h00; mem['h779E]=8'h00; mem['h779F]=8'h00;
    mem['h77A0]=8'h00; mem['h77A1]=8'h00; mem['h77A2]=8'h00; mem['h77A3]=8'h00;
    mem['h77A4]=8'h00; mem['h77A5]=8'h00; mem['h77A6]=8'h00; mem['h77A7]=8'h00;
    mem['h77A8]=8'h00; mem['h77A9]=8'h00; mem['h77AA]=8'h00; mem['h77AB]=8'h00;
    mem['h77AC]=8'h00; mem['h77AD]=8'h00; mem['h77AE]=8'h00; mem['h77AF]=8'h00;
    mem['h77B0]=8'h00; mem['h77B1]=8'h00; mem['h77B2]=8'h00; mem['h77B3]=8'h00;
    mem['h77B4]=8'h00; mem['h77B5]=8'h00; mem['h77B6]=8'h00; mem['h77B7]=8'h00;
    mem['h77B8]=8'h00; mem['h77B9]=8'h00; mem['h77BA]=8'h00; mem['h77BB]=8'h00;
    mem['h77BC]=8'h00; mem['h77BD]=8'h00; mem['h77BE]=8'h00; mem['h77BF]=8'h00;
    mem['h77C0]=8'h00; mem['h77C1]=8'h00; mem['h77C2]=8'h00; mem['h77C3]=8'h00;
    mem['h77C4]=8'h00; mem['h77C5]=8'h00; mem['h77C6]=8'h00; mem['h77C7]=8'h00;
    mem['h77C8]=8'h00; mem['h77C9]=8'h00; mem['h77CA]=8'h00; mem['h77CB]=8'h00;
    mem['h77CC]=8'h00; mem['h77CD]=8'h00; mem['h77CE]=8'h00; mem['h77CF]=8'h00;
    mem['h77D0]=8'h00; mem['h77D1]=8'h00; mem['h77D2]=8'h00; mem['h77D3]=8'h00;
    mem['h77D4]=8'h00; mem['h77D5]=8'h00; mem['h77D6]=8'h00; mem['h77D7]=8'h00;
    mem['h77D8]=8'h00; mem['h77D9]=8'h00; mem['h77DA]=8'h00; mem['h77DB]=8'h00;
    mem['h77DC]=8'h00; mem['h77DD]=8'h00; mem['h77DE]=8'h00; mem['h77DF]=8'h00;
    mem['h77E0]=8'h00; mem['h77E1]=8'h00; mem['h77E2]=8'h00; mem['h77E3]=8'h00;
    mem['h77E4]=8'h00; mem['h77E5]=8'h00; mem['h77E6]=8'h00; mem['h77E7]=8'h00;
    mem['h77E8]=8'h00; mem['h77E9]=8'h00; mem['h77EA]=8'h00; mem['h77EB]=8'h00;
    mem['h77EC]=8'h00; mem['h77ED]=8'h00; mem['h77EE]=8'h00; mem['h77EF]=8'h00;
    mem['h77F0]=8'h00; mem['h77F1]=8'h00; mem['h77F2]=8'h00; mem['h77F3]=8'h00;
    mem['h77F4]=8'h00; mem['h77F5]=8'h00; mem['h77F6]=8'h00; mem['h77F7]=8'h00;
    mem['h77F8]=8'h00; mem['h77F9]=8'h00; mem['h77FA]=8'h00; mem['h77FB]=8'h00;
    mem['h77FC]=8'h00; mem['h77FD]=8'h00; mem['h77FE]=8'h00; mem['h77FF]=8'h00;
    mem['h7800]=8'h00; mem['h7801]=8'h00; mem['h7802]=8'h00; mem['h7803]=8'h00;
    mem['h7804]=8'h00; mem['h7805]=8'h00; mem['h7806]=8'h00; mem['h7807]=8'h00;
    mem['h7808]=8'h00; mem['h7809]=8'h00; mem['h780A]=8'h00; mem['h780B]=8'h00;
    mem['h780C]=8'h00; mem['h780D]=8'h00; mem['h780E]=8'h00; mem['h780F]=8'h00;
    mem['h7810]=8'h00; mem['h7811]=8'h00; mem['h7812]=8'h00; mem['h7813]=8'h00;
    mem['h7814]=8'h00; mem['h7815]=8'h00; mem['h7816]=8'h00; mem['h7817]=8'h00;
    mem['h7818]=8'h00; mem['h7819]=8'h00; mem['h781A]=8'h00; mem['h781B]=8'h00;
    mem['h781C]=8'h00; mem['h781D]=8'h00; mem['h781E]=8'h00; mem['h781F]=8'h00;
    mem['h7820]=8'h00; mem['h7821]=8'h00; mem['h7822]=8'h00; mem['h7823]=8'h00;
    mem['h7824]=8'h00; mem['h7825]=8'h00; mem['h7826]=8'h00; mem['h7827]=8'h00;
    mem['h7828]=8'h00; mem['h7829]=8'h00; mem['h782A]=8'h00; mem['h782B]=8'h00;
    mem['h782C]=8'h00; mem['h782D]=8'h00; mem['h782E]=8'h00; mem['h782F]=8'h00;
    mem['h7830]=8'h00; mem['h7831]=8'h00; mem['h7832]=8'h00; mem['h7833]=8'h00;
    mem['h7834]=8'h00; mem['h7835]=8'h00; mem['h7836]=8'h00; mem['h7837]=8'h00;
    mem['h7838]=8'h00; mem['h7839]=8'h00; mem['h783A]=8'h00; mem['h783B]=8'h00;
    mem['h783C]=8'h00; mem['h783D]=8'h00; mem['h783E]=8'h00; mem['h783F]=8'h00;
    mem['h7840]=8'h00; mem['h7841]=8'h00; mem['h7842]=8'h00; mem['h7843]=8'h00;
    mem['h7844]=8'h00; mem['h7845]=8'h00; mem['h7846]=8'h00; mem['h7847]=8'h00;
    mem['h7848]=8'h00; mem['h7849]=8'h00; mem['h784A]=8'h00; mem['h784B]=8'h00;
    mem['h784C]=8'h00; mem['h784D]=8'h00; mem['h784E]=8'h00; mem['h784F]=8'h00;
    mem['h7850]=8'h00; mem['h7851]=8'h00; mem['h7852]=8'h00; mem['h7853]=8'h00;
    mem['h7854]=8'h00; mem['h7855]=8'h00; mem['h7856]=8'h00; mem['h7857]=8'h00;
    mem['h7858]=8'h00; mem['h7859]=8'h00; mem['h785A]=8'h00; mem['h785B]=8'h00;
    mem['h785C]=8'h00; mem['h785D]=8'h00; mem['h785E]=8'h00; mem['h785F]=8'h00;
    mem['h7860]=8'h00; mem['h7861]=8'h00; mem['h7862]=8'h00; mem['h7863]=8'h00;
    mem['h7864]=8'h00; mem['h7865]=8'h00; mem['h7866]=8'h00; mem['h7867]=8'h00;
    mem['h7868]=8'h00; mem['h7869]=8'h00; mem['h786A]=8'h00; mem['h786B]=8'h00;
    mem['h786C]=8'h00; mem['h786D]=8'h00; mem['h786E]=8'h00; mem['h786F]=8'h00;
    mem['h7870]=8'h00; mem['h7871]=8'h00; mem['h7872]=8'h00; mem['h7873]=8'h00;
    mem['h7874]=8'h00; mem['h7875]=8'h00; mem['h7876]=8'h00; mem['h7877]=8'h00;
    mem['h7878]=8'h00; mem['h7879]=8'h00; mem['h787A]=8'h00; mem['h787B]=8'h00;
    mem['h787C]=8'h00; mem['h787D]=8'h00; mem['h787E]=8'h00; mem['h787F]=8'h00;
    mem['h7880]=8'h00; mem['h7881]=8'h00; mem['h7882]=8'h00; mem['h7883]=8'h00;
    mem['h7884]=8'h00; mem['h7885]=8'h00; mem['h7886]=8'h00; mem['h7887]=8'h00;
    mem['h7888]=8'h00; mem['h7889]=8'h00; mem['h788A]=8'h00; mem['h788B]=8'h00;
    mem['h788C]=8'h00; mem['h788D]=8'h00; mem['h788E]=8'h00; mem['h788F]=8'h00;
    mem['h7890]=8'h00; mem['h7891]=8'h00; mem['h7892]=8'h00; mem['h7893]=8'h00;
    mem['h7894]=8'h00; mem['h7895]=8'h00; mem['h7896]=8'h00; mem['h7897]=8'h00;
    mem['h7898]=8'h00; mem['h7899]=8'h00; mem['h789A]=8'h00; mem['h789B]=8'h00;
    mem['h789C]=8'h00; mem['h789D]=8'h00; mem['h789E]=8'h00; mem['h789F]=8'h00;
    mem['h78A0]=8'h00; mem['h78A1]=8'h00; mem['h78A2]=8'h00; mem['h78A3]=8'h00;
    mem['h78A4]=8'h00; mem['h78A5]=8'h00; mem['h78A6]=8'h00; mem['h78A7]=8'h00;
    mem['h78A8]=8'h00; mem['h78A9]=8'h00; mem['h78AA]=8'h00; mem['h78AB]=8'h00;
    mem['h78AC]=8'h00; mem['h78AD]=8'h00; mem['h78AE]=8'h00; mem['h78AF]=8'h00;
    mem['h78B0]=8'h00; mem['h78B1]=8'h00; mem['h78B2]=8'h00; mem['h78B3]=8'h00;
    mem['h78B4]=8'h00; mem['h78B5]=8'h00; mem['h78B6]=8'h00; mem['h78B7]=8'h00;
    mem['h78B8]=8'h00; mem['h78B9]=8'h00; mem['h78BA]=8'h00; mem['h78BB]=8'h00;
    mem['h78BC]=8'h00; mem['h78BD]=8'h00; mem['h78BE]=8'h00; mem['h78BF]=8'h00;
    mem['h78C0]=8'h00; mem['h78C1]=8'h00; mem['h78C2]=8'h00; mem['h78C3]=8'h00;
    mem['h78C4]=8'h00; mem['h78C5]=8'h00; mem['h78C6]=8'h00; mem['h78C7]=8'h00;
    mem['h78C8]=8'h00; mem['h78C9]=8'h00; mem['h78CA]=8'h00; mem['h78CB]=8'h00;
    mem['h78CC]=8'h00; mem['h78CD]=8'h00; mem['h78CE]=8'h00; mem['h78CF]=8'h00;
    mem['h78D0]=8'h00; mem['h78D1]=8'h00; mem['h78D2]=8'h00; mem['h78D3]=8'h00;
    mem['h78D4]=8'h00; mem['h78D5]=8'h00; mem['h78D6]=8'h00; mem['h78D7]=8'h00;
    mem['h78D8]=8'h00; mem['h78D9]=8'h00; mem['h78DA]=8'h00; mem['h78DB]=8'h00;
    mem['h78DC]=8'h00; mem['h78DD]=8'h00; mem['h78DE]=8'h00; mem['h78DF]=8'h00;
    mem['h78E0]=8'h00; mem['h78E1]=8'h00; mem['h78E2]=8'h00; mem['h78E3]=8'h00;
    mem['h78E4]=8'h00; mem['h78E5]=8'h00; mem['h78E6]=8'h00; mem['h78E7]=8'h00;
    mem['h78E8]=8'h00; mem['h78E9]=8'h00; mem['h78EA]=8'h00; mem['h78EB]=8'h00;
    mem['h78EC]=8'h00; mem['h78ED]=8'h00; mem['h78EE]=8'h00; mem['h78EF]=8'h00;
    mem['h78F0]=8'h00; mem['h78F1]=8'h00; mem['h78F2]=8'h00; mem['h78F3]=8'h00;
    mem['h78F4]=8'h00; mem['h78F5]=8'h00; mem['h78F6]=8'h00; mem['h78F7]=8'h00;
    mem['h78F8]=8'h00; mem['h78F9]=8'h00; mem['h78FA]=8'h00; mem['h78FB]=8'h00;
    mem['h78FC]=8'h00; mem['h78FD]=8'h00; mem['h78FE]=8'h00; mem['h78FF]=8'h00;
    mem['h7900]=8'h00; mem['h7901]=8'h00; mem['h7902]=8'h00; mem['h7903]=8'h00;
    mem['h7904]=8'h00; mem['h7905]=8'h00; mem['h7906]=8'h00; mem['h7907]=8'h00;
    mem['h7908]=8'h00; mem['h7909]=8'h00; mem['h790A]=8'h00; mem['h790B]=8'h00;
    mem['h790C]=8'h00; mem['h790D]=8'h00; mem['h790E]=8'h00; mem['h790F]=8'h00;
    mem['h7910]=8'h00; mem['h7911]=8'h00; mem['h7912]=8'h00; mem['h7913]=8'h00;
    mem['h7914]=8'h00; mem['h7915]=8'h00; mem['h7916]=8'h00; mem['h7917]=8'h00;
    mem['h7918]=8'h00; mem['h7919]=8'h00; mem['h791A]=8'h00; mem['h791B]=8'h00;
    mem['h791C]=8'h00; mem['h791D]=8'h00; mem['h791E]=8'h00; mem['h791F]=8'h00;
    mem['h7920]=8'h00; mem['h7921]=8'h00; mem['h7922]=8'h00; mem['h7923]=8'h00;
    mem['h7924]=8'h00; mem['h7925]=8'h00; mem['h7926]=8'h00; mem['h7927]=8'h00;
    mem['h7928]=8'h00; mem['h7929]=8'h00; mem['h792A]=8'h00; mem['h792B]=8'h00;
    mem['h792C]=8'h00; mem['h792D]=8'h00; mem['h792E]=8'h00; mem['h792F]=8'h00;
    mem['h7930]=8'h00; mem['h7931]=8'h00; mem['h7932]=8'h00; mem['h7933]=8'h00;
    mem['h7934]=8'h00; mem['h7935]=8'h00; mem['h7936]=8'h00; mem['h7937]=8'h00;
    mem['h7938]=8'h00; mem['h7939]=8'h00; mem['h793A]=8'h00; mem['h793B]=8'h00;
    mem['h793C]=8'h00; mem['h793D]=8'h00; mem['h793E]=8'h00; mem['h793F]=8'h00;
    mem['h7940]=8'h00; mem['h7941]=8'h00; mem['h7942]=8'h00; mem['h7943]=8'h00;
    mem['h7944]=8'h00; mem['h7945]=8'h00; mem['h7946]=8'h00; mem['h7947]=8'h00;
    mem['h7948]=8'h00; mem['h7949]=8'h00; mem['h794A]=8'h00; mem['h794B]=8'h00;
    mem['h794C]=8'h00; mem['h794D]=8'h00; mem['h794E]=8'h00; mem['h794F]=8'h00;
    mem['h7950]=8'h00; mem['h7951]=8'h00; mem['h7952]=8'h00; mem['h7953]=8'h00;
    mem['h7954]=8'h00; mem['h7955]=8'h00; mem['h7956]=8'h00; mem['h7957]=8'h00;
    mem['h7958]=8'h00; mem['h7959]=8'h00; mem['h795A]=8'h00; mem['h795B]=8'h00;
    mem['h795C]=8'h00; mem['h795D]=8'h00; mem['h795E]=8'h00; mem['h795F]=8'h00;
    mem['h7960]=8'h00; mem['h7961]=8'h00; mem['h7962]=8'h00; mem['h7963]=8'h00;
    mem['h7964]=8'h00; mem['h7965]=8'h00; mem['h7966]=8'h00; mem['h7967]=8'h00;
    mem['h7968]=8'h00; mem['h7969]=8'h00; mem['h796A]=8'h00; mem['h796B]=8'h00;
    mem['h796C]=8'h00; mem['h796D]=8'h00; mem['h796E]=8'h00; mem['h796F]=8'h00;
    mem['h7970]=8'h00; mem['h7971]=8'h00; mem['h7972]=8'h00; mem['h7973]=8'h00;
    mem['h7974]=8'h00; mem['h7975]=8'h00; mem['h7976]=8'h00; mem['h7977]=8'h00;
    mem['h7978]=8'h00; mem['h7979]=8'h00; mem['h797A]=8'h00; mem['h797B]=8'h00;
    mem['h797C]=8'h00; mem['h797D]=8'h00; mem['h797E]=8'h00; mem['h797F]=8'h00;
    mem['h7980]=8'h00; mem['h7981]=8'h00; mem['h7982]=8'h00; mem['h7983]=8'h00;
    mem['h7984]=8'h00; mem['h7985]=8'h00; mem['h7986]=8'h00; mem['h7987]=8'h00;
    mem['h7988]=8'h00; mem['h7989]=8'h00; mem['h798A]=8'h00; mem['h798B]=8'h00;
    mem['h798C]=8'h00; mem['h798D]=8'h00; mem['h798E]=8'h00; mem['h798F]=8'h00;
    mem['h7990]=8'h00; mem['h7991]=8'h00; mem['h7992]=8'h00; mem['h7993]=8'h00;
    mem['h7994]=8'h00; mem['h7995]=8'h00; mem['h7996]=8'h00; mem['h7997]=8'h00;
    mem['h7998]=8'h00; mem['h7999]=8'h00; mem['h799A]=8'h00; mem['h799B]=8'h00;
    mem['h799C]=8'h00; mem['h799D]=8'h00; mem['h799E]=8'h00; mem['h799F]=8'h00;
    mem['h79A0]=8'h00; mem['h79A1]=8'h00; mem['h79A2]=8'h00; mem['h79A3]=8'h00;
    mem['h79A4]=8'h00; mem['h79A5]=8'h00; mem['h79A6]=8'h00; mem['h79A7]=8'h00;
    mem['h79A8]=8'h00; mem['h79A9]=8'h00; mem['h79AA]=8'h00; mem['h79AB]=8'h00;
    mem['h79AC]=8'h00; mem['h79AD]=8'h00; mem['h79AE]=8'h00; mem['h79AF]=8'h00;
    mem['h79B0]=8'h00; mem['h79B1]=8'h00; mem['h79B2]=8'h00; mem['h79B3]=8'h00;
    mem['h79B4]=8'h00; mem['h79B5]=8'h00; mem['h79B6]=8'h00; mem['h79B7]=8'h00;
    mem['h79B8]=8'h00; mem['h79B9]=8'h00; mem['h79BA]=8'h00; mem['h79BB]=8'h00;
    mem['h79BC]=8'h00; mem['h79BD]=8'h00; mem['h79BE]=8'h00; mem['h79BF]=8'h00;
    mem['h79C0]=8'h00; mem['h79C1]=8'h00; mem['h79C2]=8'h00; mem['h79C3]=8'h00;
    mem['h79C4]=8'h00; mem['h79C5]=8'h00; mem['h79C6]=8'h00; mem['h79C7]=8'h00;
    mem['h79C8]=8'h00; mem['h79C9]=8'h00; mem['h79CA]=8'h00; mem['h79CB]=8'h00;
    mem['h79CC]=8'h00; mem['h79CD]=8'h00; mem['h79CE]=8'h00; mem['h79CF]=8'h00;
    mem['h79D0]=8'h00; mem['h79D1]=8'h00; mem['h79D2]=8'h00; mem['h79D3]=8'h00;
    mem['h79D4]=8'h00; mem['h79D5]=8'h00; mem['h79D6]=8'h00; mem['h79D7]=8'h00;
    mem['h79D8]=8'h00; mem['h79D9]=8'h00; mem['h79DA]=8'h00; mem['h79DB]=8'h00;
    mem['h79DC]=8'h00; mem['h79DD]=8'h00; mem['h79DE]=8'h00; mem['h79DF]=8'h00;
    mem['h79E0]=8'h00; mem['h79E1]=8'h00; mem['h79E2]=8'h00; mem['h79E3]=8'h00;
    mem['h79E4]=8'h00; mem['h79E5]=8'h00; mem['h79E6]=8'h00; mem['h79E7]=8'h00;
    mem['h79E8]=8'h00; mem['h79E9]=8'h00; mem['h79EA]=8'h00; mem['h79EB]=8'h00;
    mem['h79EC]=8'h00; mem['h79ED]=8'h00; mem['h79EE]=8'h00; mem['h79EF]=8'h00;
    mem['h79F0]=8'h00; mem['h79F1]=8'h00; mem['h79F2]=8'h00; mem['h79F3]=8'h00;
    mem['h79F4]=8'h00; mem['h79F5]=8'h00; mem['h79F6]=8'h00; mem['h79F7]=8'h00;
    mem['h79F8]=8'h00; mem['h79F9]=8'h00; mem['h79FA]=8'h00; mem['h79FB]=8'h00;
    mem['h79FC]=8'h00; mem['h79FD]=8'h00; mem['h79FE]=8'h00; mem['h79FF]=8'h00;
    mem['h7A00]=8'h00; mem['h7A01]=8'h00; mem['h7A02]=8'h00; mem['h7A03]=8'h00;
    mem['h7A04]=8'h00; mem['h7A05]=8'h00; mem['h7A06]=8'h00; mem['h7A07]=8'h00;
    mem['h7A08]=8'h00; mem['h7A09]=8'h00; mem['h7A0A]=8'h00; mem['h7A0B]=8'h00;
    mem['h7A0C]=8'h00; mem['h7A0D]=8'h00; mem['h7A0E]=8'h00; mem['h7A0F]=8'h00;
    mem['h7A10]=8'h00; mem['h7A11]=8'h00; mem['h7A12]=8'h00; mem['h7A13]=8'h00;
    mem['h7A14]=8'h00; mem['h7A15]=8'h00; mem['h7A16]=8'h00; mem['h7A17]=8'h00;
    mem['h7A18]=8'h00; mem['h7A19]=8'h00; mem['h7A1A]=8'h00; mem['h7A1B]=8'h00;
    mem['h7A1C]=8'h00; mem['h7A1D]=8'h00; mem['h7A1E]=8'h00; mem['h7A1F]=8'h00;
    mem['h7A20]=8'h00; mem['h7A21]=8'h00; mem['h7A22]=8'h00; mem['h7A23]=8'h00;
    mem['h7A24]=8'h00; mem['h7A25]=8'h00; mem['h7A26]=8'h00; mem['h7A27]=8'h00;
    mem['h7A28]=8'h00; mem['h7A29]=8'h00; mem['h7A2A]=8'h00; mem['h7A2B]=8'h00;
    mem['h7A2C]=8'h00; mem['h7A2D]=8'h00; mem['h7A2E]=8'h00; mem['h7A2F]=8'h00;
    mem['h7A30]=8'h00; mem['h7A31]=8'h00; mem['h7A32]=8'h00; mem['h7A33]=8'h00;
    mem['h7A34]=8'h00; mem['h7A35]=8'h00; mem['h7A36]=8'h00; mem['h7A37]=8'h00;
    mem['h7A38]=8'h00; mem['h7A39]=8'h00; mem['h7A3A]=8'h00; mem['h7A3B]=8'h00;
    mem['h7A3C]=8'h00; mem['h7A3D]=8'h00; mem['h7A3E]=8'h00; mem['h7A3F]=8'h00;
    mem['h7A40]=8'h00; mem['h7A41]=8'h00; mem['h7A42]=8'h00; mem['h7A43]=8'h00;
    mem['h7A44]=8'h00; mem['h7A45]=8'h00; mem['h7A46]=8'h00; mem['h7A47]=8'h00;
    mem['h7A48]=8'h00; mem['h7A49]=8'h00; mem['h7A4A]=8'h00; mem['h7A4B]=8'h00;
    mem['h7A4C]=8'h00; mem['h7A4D]=8'h00; mem['h7A4E]=8'h00; mem['h7A4F]=8'h00;
    mem['h7A50]=8'h00; mem['h7A51]=8'h00; mem['h7A52]=8'h00; mem['h7A53]=8'h00;
    mem['h7A54]=8'h00; mem['h7A55]=8'h00; mem['h7A56]=8'h00; mem['h7A57]=8'h00;
    mem['h7A58]=8'h00; mem['h7A59]=8'h00; mem['h7A5A]=8'h00; mem['h7A5B]=8'h00;
    mem['h7A5C]=8'h00; mem['h7A5D]=8'h00; mem['h7A5E]=8'h00; mem['h7A5F]=8'h00;
    mem['h7A60]=8'h00; mem['h7A61]=8'h00; mem['h7A62]=8'h00; mem['h7A63]=8'h00;
    mem['h7A64]=8'h00; mem['h7A65]=8'h00; mem['h7A66]=8'h00; mem['h7A67]=8'h00;
    mem['h7A68]=8'h00; mem['h7A69]=8'h00; mem['h7A6A]=8'h00; mem['h7A6B]=8'h00;
    mem['h7A6C]=8'h00; mem['h7A6D]=8'h00; mem['h7A6E]=8'h00; mem['h7A6F]=8'h00;
    mem['h7A70]=8'h00; mem['h7A71]=8'h00; mem['h7A72]=8'h00; mem['h7A73]=8'h00;
    mem['h7A74]=8'h00; mem['h7A75]=8'h00; mem['h7A76]=8'h00; mem['h7A77]=8'h00;
    mem['h7A78]=8'h00; mem['h7A79]=8'h00; mem['h7A7A]=8'h00; mem['h7A7B]=8'h00;
    mem['h7A7C]=8'h00; mem['h7A7D]=8'h00; mem['h7A7E]=8'h00; mem['h7A7F]=8'h00;
    mem['h7A80]=8'h00; mem['h7A81]=8'h00; mem['h7A82]=8'h00; mem['h7A83]=8'h00;
    mem['h7A84]=8'h00; mem['h7A85]=8'h00; mem['h7A86]=8'h00; mem['h7A87]=8'h00;
    mem['h7A88]=8'h00; mem['h7A89]=8'h00; mem['h7A8A]=8'h00; mem['h7A8B]=8'h00;
    mem['h7A8C]=8'h00; mem['h7A8D]=8'h00; mem['h7A8E]=8'h00; mem['h7A8F]=8'h00;
    mem['h7A90]=8'h00; mem['h7A91]=8'h00; mem['h7A92]=8'h00; mem['h7A93]=8'h00;
    mem['h7A94]=8'h00; mem['h7A95]=8'h00; mem['h7A96]=8'h00; mem['h7A97]=8'h00;
    mem['h7A98]=8'h00; mem['h7A99]=8'h00; mem['h7A9A]=8'h00; mem['h7A9B]=8'h00;
    mem['h7A9C]=8'h00; mem['h7A9D]=8'h00; mem['h7A9E]=8'h00; mem['h7A9F]=8'h00;
    mem['h7AA0]=8'h00; mem['h7AA1]=8'h00; mem['h7AA2]=8'h00; mem['h7AA3]=8'h00;
    mem['h7AA4]=8'h00; mem['h7AA5]=8'h00; mem['h7AA6]=8'h00; mem['h7AA7]=8'h00;
    mem['h7AA8]=8'h00; mem['h7AA9]=8'h00; mem['h7AAA]=8'h00; mem['h7AAB]=8'h00;
    mem['h7AAC]=8'h00; mem['h7AAD]=8'h00; mem['h7AAE]=8'h00; mem['h7AAF]=8'h00;
    mem['h7AB0]=8'h00; mem['h7AB1]=8'h00; mem['h7AB2]=8'h00; mem['h7AB3]=8'h00;
    mem['h7AB4]=8'h00; mem['h7AB5]=8'h00; mem['h7AB6]=8'h00; mem['h7AB7]=8'h00;
    mem['h7AB8]=8'h00; mem['h7AB9]=8'h00; mem['h7ABA]=8'h00; mem['h7ABB]=8'h00;
    mem['h7ABC]=8'h00; mem['h7ABD]=8'h00; mem['h7ABE]=8'h00; mem['h7ABF]=8'h00;
    mem['h7AC0]=8'h00; mem['h7AC1]=8'h00; mem['h7AC2]=8'h00; mem['h7AC3]=8'h00;
    mem['h7AC4]=8'h00; mem['h7AC5]=8'h00; mem['h7AC6]=8'h00; mem['h7AC7]=8'h00;
    mem['h7AC8]=8'h00; mem['h7AC9]=8'h00; mem['h7ACA]=8'h00; mem['h7ACB]=8'h00;
    mem['h7ACC]=8'h00; mem['h7ACD]=8'h00; mem['h7ACE]=8'h00; mem['h7ACF]=8'h00;
    mem['h7AD0]=8'h00; mem['h7AD1]=8'h00; mem['h7AD2]=8'h00; mem['h7AD3]=8'h00;
    mem['h7AD4]=8'h00; mem['h7AD5]=8'h00; mem['h7AD6]=8'h00; mem['h7AD7]=8'h00;
    mem['h7AD8]=8'h00; mem['h7AD9]=8'h00; mem['h7ADA]=8'h00; mem['h7ADB]=8'h00;
    mem['h7ADC]=8'h00; mem['h7ADD]=8'h00; mem['h7ADE]=8'h00; mem['h7ADF]=8'h00;
    mem['h7AE0]=8'h00; mem['h7AE1]=8'h00; mem['h7AE2]=8'h00; mem['h7AE3]=8'h00;
    mem['h7AE4]=8'h00; mem['h7AE5]=8'h00; mem['h7AE6]=8'h00; mem['h7AE7]=8'h00;
    mem['h7AE8]=8'h00; mem['h7AE9]=8'h00; mem['h7AEA]=8'h00; mem['h7AEB]=8'h00;
    mem['h7AEC]=8'h00; mem['h7AED]=8'h00; mem['h7AEE]=8'h00; mem['h7AEF]=8'h00;
    mem['h7AF0]=8'h00; mem['h7AF1]=8'h00; mem['h7AF2]=8'h00; mem['h7AF3]=8'h00;
    mem['h7AF4]=8'h00; mem['h7AF5]=8'h00; mem['h7AF6]=8'h00; mem['h7AF7]=8'h00;
    mem['h7AF8]=8'h00; mem['h7AF9]=8'h00; mem['h7AFA]=8'h00; mem['h7AFB]=8'h00;
    mem['h7AFC]=8'h00; mem['h7AFD]=8'h00; mem['h7AFE]=8'h00; mem['h7AFF]=8'h00;
    mem['h7B00]=8'h00; mem['h7B01]=8'h00; mem['h7B02]=8'h00; mem['h7B03]=8'h00;
    mem['h7B04]=8'h00; mem['h7B05]=8'h00; mem['h7B06]=8'h00; mem['h7B07]=8'h00;
    mem['h7B08]=8'h00; mem['h7B09]=8'h00; mem['h7B0A]=8'h00; mem['h7B0B]=8'h00;
    mem['h7B0C]=8'h00; mem['h7B0D]=8'h00; mem['h7B0E]=8'h00; mem['h7B0F]=8'h00;
    mem['h7B10]=8'h00; mem['h7B11]=8'h00; mem['h7B12]=8'h00; mem['h7B13]=8'h00;
    mem['h7B14]=8'h00; mem['h7B15]=8'h00; mem['h7B16]=8'h00; mem['h7B17]=8'h00;
    mem['h7B18]=8'h00; mem['h7B19]=8'h00; mem['h7B1A]=8'h00; mem['h7B1B]=8'h00;
    mem['h7B1C]=8'h00; mem['h7B1D]=8'h00; mem['h7B1E]=8'h00; mem['h7B1F]=8'h00;
    mem['h7B20]=8'h00; mem['h7B21]=8'h00; mem['h7B22]=8'h00; mem['h7B23]=8'h00;
    mem['h7B24]=8'h00; mem['h7B25]=8'h00; mem['h7B26]=8'h00; mem['h7B27]=8'h00;
    mem['h7B28]=8'h00; mem['h7B29]=8'h00; mem['h7B2A]=8'h00; mem['h7B2B]=8'h00;
    mem['h7B2C]=8'h00; mem['h7B2D]=8'h00; mem['h7B2E]=8'h00; mem['h7B2F]=8'h00;
    mem['h7B30]=8'h00; mem['h7B31]=8'h00; mem['h7B32]=8'h00; mem['h7B33]=8'h00;
    mem['h7B34]=8'h00; mem['h7B35]=8'h00; mem['h7B36]=8'h00; mem['h7B37]=8'h00;
    mem['h7B38]=8'h00; mem['h7B39]=8'h00; mem['h7B3A]=8'h00; mem['h7B3B]=8'h00;
    mem['h7B3C]=8'h00; mem['h7B3D]=8'h00; mem['h7B3E]=8'h00; mem['h7B3F]=8'h00;
    mem['h7B40]=8'h00; mem['h7B41]=8'h00; mem['h7B42]=8'h00; mem['h7B43]=8'h00;
    mem['h7B44]=8'h00; mem['h7B45]=8'h00; mem['h7B46]=8'h00; mem['h7B47]=8'h00;
    mem['h7B48]=8'h00; mem['h7B49]=8'h00; mem['h7B4A]=8'h00; mem['h7B4B]=8'h00;
    mem['h7B4C]=8'h00; mem['h7B4D]=8'h00; mem['h7B4E]=8'h00; mem['h7B4F]=8'h00;
    mem['h7B50]=8'h00; mem['h7B51]=8'h00; mem['h7B52]=8'h00; mem['h7B53]=8'h00;
    mem['h7B54]=8'h00; mem['h7B55]=8'h00; mem['h7B56]=8'h00; mem['h7B57]=8'h00;
    mem['h7B58]=8'h00; mem['h7B59]=8'h00; mem['h7B5A]=8'h00; mem['h7B5B]=8'h00;
    mem['h7B5C]=8'h00; mem['h7B5D]=8'h00; mem['h7B5E]=8'h00; mem['h7B5F]=8'h00;
    mem['h7B60]=8'h00; mem['h7B61]=8'h00; mem['h7B62]=8'h00; mem['h7B63]=8'h00;
    mem['h7B64]=8'h00; mem['h7B65]=8'h00; mem['h7B66]=8'h00; mem['h7B67]=8'h00;
    mem['h7B68]=8'h00; mem['h7B69]=8'h00; mem['h7B6A]=8'h00; mem['h7B6B]=8'h00;
    mem['h7B6C]=8'h00; mem['h7B6D]=8'h00; mem['h7B6E]=8'h00; mem['h7B6F]=8'h00;
    mem['h7B70]=8'h00; mem['h7B71]=8'h00; mem['h7B72]=8'h00; mem['h7B73]=8'h00;
    mem['h7B74]=8'h00; mem['h7B75]=8'h00; mem['h7B76]=8'h00; mem['h7B77]=8'h00;
    mem['h7B78]=8'h00; mem['h7B79]=8'h00; mem['h7B7A]=8'h00; mem['h7B7B]=8'h00;
    mem['h7B7C]=8'h00; mem['h7B7D]=8'h00; mem['h7B7E]=8'h00; mem['h7B7F]=8'h00;
    mem['h7B80]=8'h00; mem['h7B81]=8'h00; mem['h7B82]=8'h00; mem['h7B83]=8'h00;
    mem['h7B84]=8'h00; mem['h7B85]=8'h00; mem['h7B86]=8'h00; mem['h7B87]=8'h00;
    mem['h7B88]=8'h00; mem['h7B89]=8'h00; mem['h7B8A]=8'h00; mem['h7B8B]=8'h00;
    mem['h7B8C]=8'h00; mem['h7B8D]=8'h00; mem['h7B8E]=8'h00; mem['h7B8F]=8'h00;
    mem['h7B90]=8'h00; mem['h7B91]=8'h00; mem['h7B92]=8'h00; mem['h7B93]=8'h00;
    mem['h7B94]=8'h00; mem['h7B95]=8'h00; mem['h7B96]=8'h00; mem['h7B97]=8'h00;
    mem['h7B98]=8'h00; mem['h7B99]=8'h00; mem['h7B9A]=8'h00; mem['h7B9B]=8'h00;
    mem['h7B9C]=8'h00; mem['h7B9D]=8'h00; mem['h7B9E]=8'h00; mem['h7B9F]=8'h00;
    mem['h7BA0]=8'h00; mem['h7BA1]=8'h00; mem['h7BA2]=8'h00; mem['h7BA3]=8'h00;
    mem['h7BA4]=8'h00; mem['h7BA5]=8'h00; mem['h7BA6]=8'h00; mem['h7BA7]=8'h00;
    mem['h7BA8]=8'h00; mem['h7BA9]=8'h00; mem['h7BAA]=8'h00; mem['h7BAB]=8'h00;
    mem['h7BAC]=8'h00; mem['h7BAD]=8'h00; mem['h7BAE]=8'h00; mem['h7BAF]=8'h00;
    mem['h7BB0]=8'h00; mem['h7BB1]=8'h00; mem['h7BB2]=8'h00; mem['h7BB3]=8'h00;
    mem['h7BB4]=8'h00; mem['h7BB5]=8'h00; mem['h7BB6]=8'h00; mem['h7BB7]=8'h00;
    mem['h7BB8]=8'h00; mem['h7BB9]=8'h00; mem['h7BBA]=8'h00; mem['h7BBB]=8'h00;
    mem['h7BBC]=8'h00; mem['h7BBD]=8'h00; mem['h7BBE]=8'h00; mem['h7BBF]=8'h00;
    mem['h7BC0]=8'h00; mem['h7BC1]=8'h00; mem['h7BC2]=8'h00; mem['h7BC3]=8'h00;
    mem['h7BC4]=8'h00; mem['h7BC5]=8'h00; mem['h7BC6]=8'h00; mem['h7BC7]=8'h00;
    mem['h7BC8]=8'h00; mem['h7BC9]=8'h00; mem['h7BCA]=8'h00; mem['h7BCB]=8'h00;
    mem['h7BCC]=8'h00; mem['h7BCD]=8'h00; mem['h7BCE]=8'h00; mem['h7BCF]=8'h00;
    mem['h7BD0]=8'h00; mem['h7BD1]=8'h00; mem['h7BD2]=8'h00; mem['h7BD3]=8'h00;
    mem['h7BD4]=8'h00; mem['h7BD5]=8'h00; mem['h7BD6]=8'h00; mem['h7BD7]=8'h00;
    mem['h7BD8]=8'h00; mem['h7BD9]=8'h00; mem['h7BDA]=8'h00; mem['h7BDB]=8'h00;
    mem['h7BDC]=8'h00; mem['h7BDD]=8'h00; mem['h7BDE]=8'h00; mem['h7BDF]=8'h00;
    mem['h7BE0]=8'h00; mem['h7BE1]=8'h00; mem['h7BE2]=8'h00; mem['h7BE3]=8'h00;
    mem['h7BE4]=8'h00; mem['h7BE5]=8'h00; mem['h7BE6]=8'h00; mem['h7BE7]=8'h00;
    mem['h7BE8]=8'h00; mem['h7BE9]=8'h00; mem['h7BEA]=8'h00; mem['h7BEB]=8'h00;
    mem['h7BEC]=8'h00; mem['h7BED]=8'h00; mem['h7BEE]=8'h00; mem['h7BEF]=8'h00;
    mem['h7BF0]=8'h00; mem['h7BF1]=8'h00; mem['h7BF2]=8'h00; mem['h7BF3]=8'h00;
    mem['h7BF4]=8'h00; mem['h7BF5]=8'h00; mem['h7BF6]=8'h00; mem['h7BF7]=8'h00;
    mem['h7BF8]=8'h00; mem['h7BF9]=8'h00; mem['h7BFA]=8'h00; mem['h7BFB]=8'h00;
    mem['h7BFC]=8'h00; mem['h7BFD]=8'h00; mem['h7BFE]=8'h00; mem['h7BFF]=8'h00;
    mem['h7C00]=8'h00; mem['h7C01]=8'h00; mem['h7C02]=8'h00; mem['h7C03]=8'h00;
    mem['h7C04]=8'h00; mem['h7C05]=8'h00; mem['h7C06]=8'h00; mem['h7C07]=8'h00;
    mem['h7C08]=8'h00; mem['h7C09]=8'h00; mem['h7C0A]=8'h00; mem['h7C0B]=8'h00;
    mem['h7C0C]=8'h00; mem['h7C0D]=8'h00; mem['h7C0E]=8'h00; mem['h7C0F]=8'h00;
    mem['h7C10]=8'h00; mem['h7C11]=8'h00; mem['h7C12]=8'h00; mem['h7C13]=8'h00;
    mem['h7C14]=8'h00; mem['h7C15]=8'h00; mem['h7C16]=8'h00; mem['h7C17]=8'h00;
    mem['h7C18]=8'h00; mem['h7C19]=8'h00; mem['h7C1A]=8'h00; mem['h7C1B]=8'h00;
    mem['h7C1C]=8'h00; mem['h7C1D]=8'h00; mem['h7C1E]=8'h00; mem['h7C1F]=8'h00;
    mem['h7C20]=8'h00; mem['h7C21]=8'h00; mem['h7C22]=8'h00; mem['h7C23]=8'h00;
    mem['h7C24]=8'h00; mem['h7C25]=8'h00; mem['h7C26]=8'h00; mem['h7C27]=8'h00;
    mem['h7C28]=8'h00; mem['h7C29]=8'h00; mem['h7C2A]=8'h00; mem['h7C2B]=8'h00;
    mem['h7C2C]=8'h00; mem['h7C2D]=8'h00; mem['h7C2E]=8'h00; mem['h7C2F]=8'h00;
    mem['h7C30]=8'h00; mem['h7C31]=8'h00; mem['h7C32]=8'h00; mem['h7C33]=8'h00;
    mem['h7C34]=8'h00; mem['h7C35]=8'h00; mem['h7C36]=8'h00; mem['h7C37]=8'h00;
    mem['h7C38]=8'h00; mem['h7C39]=8'h00; mem['h7C3A]=8'h00; mem['h7C3B]=8'h00;
    mem['h7C3C]=8'h00; mem['h7C3D]=8'h00; mem['h7C3E]=8'h00; mem['h7C3F]=8'h00;
    mem['h7C40]=8'h00; mem['h7C41]=8'h00; mem['h7C42]=8'h00; mem['h7C43]=8'h00;
    mem['h7C44]=8'h00; mem['h7C45]=8'h00; mem['h7C46]=8'h00; mem['h7C47]=8'h00;
    mem['h7C48]=8'h00; mem['h7C49]=8'h00; mem['h7C4A]=8'h00; mem['h7C4B]=8'h00;
    mem['h7C4C]=8'h00; mem['h7C4D]=8'h00; mem['h7C4E]=8'h00; mem['h7C4F]=8'h00;
    mem['h7C50]=8'h00; mem['h7C51]=8'h00; mem['h7C52]=8'h00; mem['h7C53]=8'h00;
    mem['h7C54]=8'h00; mem['h7C55]=8'h00; mem['h7C56]=8'h00; mem['h7C57]=8'h00;
    mem['h7C58]=8'h00; mem['h7C59]=8'h00; mem['h7C5A]=8'h00; mem['h7C5B]=8'h00;
    mem['h7C5C]=8'h00; mem['h7C5D]=8'h00; mem['h7C5E]=8'h00; mem['h7C5F]=8'h00;
    mem['h7C60]=8'h00; mem['h7C61]=8'h00; mem['h7C62]=8'h00; mem['h7C63]=8'h00;
    mem['h7C64]=8'h00; mem['h7C65]=8'h00; mem['h7C66]=8'h00; mem['h7C67]=8'h00;
    mem['h7C68]=8'h00; mem['h7C69]=8'h00; mem['h7C6A]=8'h00; mem['h7C6B]=8'h00;
    mem['h7C6C]=8'h00; mem['h7C6D]=8'h00; mem['h7C6E]=8'h00; mem['h7C6F]=8'h00;
    mem['h7C70]=8'h00; mem['h7C71]=8'h00; mem['h7C72]=8'h00; mem['h7C73]=8'h00;
    mem['h7C74]=8'h00; mem['h7C75]=8'h00; mem['h7C76]=8'h00; mem['h7C77]=8'h00;
    mem['h7C78]=8'h00; mem['h7C79]=8'h00; mem['h7C7A]=8'h00; mem['h7C7B]=8'h00;
    mem['h7C7C]=8'h00; mem['h7C7D]=8'h00; mem['h7C7E]=8'h00; mem['h7C7F]=8'h00;
    mem['h7C80]=8'h00; mem['h7C81]=8'h00; mem['h7C82]=8'h00; mem['h7C83]=8'h00;
    mem['h7C84]=8'h00; mem['h7C85]=8'h00; mem['h7C86]=8'h00; mem['h7C87]=8'h00;
    mem['h7C88]=8'h00; mem['h7C89]=8'h00; mem['h7C8A]=8'h00; mem['h7C8B]=8'h00;
    mem['h7C8C]=8'h00; mem['h7C8D]=8'h00; mem['h7C8E]=8'h00; mem['h7C8F]=8'h00;
    mem['h7C90]=8'h00; mem['h7C91]=8'h00; mem['h7C92]=8'h00; mem['h7C93]=8'h00;
    mem['h7C94]=8'h00; mem['h7C95]=8'h00; mem['h7C96]=8'h00; mem['h7C97]=8'h00;
    mem['h7C98]=8'h00; mem['h7C99]=8'h00; mem['h7C9A]=8'h00; mem['h7C9B]=8'h00;
    mem['h7C9C]=8'h00; mem['h7C9D]=8'h00; mem['h7C9E]=8'h00; mem['h7C9F]=8'h00;
    mem['h7CA0]=8'h00; mem['h7CA1]=8'h00; mem['h7CA2]=8'h00; mem['h7CA3]=8'h00;
    mem['h7CA4]=8'h00; mem['h7CA5]=8'h00; mem['h7CA6]=8'h00; mem['h7CA7]=8'h00;
    mem['h7CA8]=8'h00; mem['h7CA9]=8'h00; mem['h7CAA]=8'h00; mem['h7CAB]=8'h00;
    mem['h7CAC]=8'h00; mem['h7CAD]=8'h00; mem['h7CAE]=8'h00; mem['h7CAF]=8'h00;
    mem['h7CB0]=8'h00; mem['h7CB1]=8'h00; mem['h7CB2]=8'h00; mem['h7CB3]=8'h00;
    mem['h7CB4]=8'h00; mem['h7CB5]=8'h00; mem['h7CB6]=8'h00; mem['h7CB7]=8'h00;
    mem['h7CB8]=8'h00; mem['h7CB9]=8'h00; mem['h7CBA]=8'h00; mem['h7CBB]=8'h00;
    mem['h7CBC]=8'h00; mem['h7CBD]=8'h00; mem['h7CBE]=8'h00; mem['h7CBF]=8'h00;
    mem['h7CC0]=8'h00; mem['h7CC1]=8'h00; mem['h7CC2]=8'h00; mem['h7CC3]=8'h00;
    mem['h7CC4]=8'h00; mem['h7CC5]=8'h00; mem['h7CC6]=8'h00; mem['h7CC7]=8'h00;
    mem['h7CC8]=8'h00; mem['h7CC9]=8'h00; mem['h7CCA]=8'h00; mem['h7CCB]=8'h00;
    mem['h7CCC]=8'h00; mem['h7CCD]=8'h00; mem['h7CCE]=8'h00; mem['h7CCF]=8'h00;
    mem['h7CD0]=8'h00; mem['h7CD1]=8'h00; mem['h7CD2]=8'h00; mem['h7CD3]=8'h00;
    mem['h7CD4]=8'h00; mem['h7CD5]=8'h00; mem['h7CD6]=8'h00; mem['h7CD7]=8'h00;
    mem['h7CD8]=8'h00; mem['h7CD9]=8'h00; mem['h7CDA]=8'h00; mem['h7CDB]=8'h00;
    mem['h7CDC]=8'h00; mem['h7CDD]=8'h00; mem['h7CDE]=8'h00; mem['h7CDF]=8'h00;
    mem['h7CE0]=8'h00; mem['h7CE1]=8'h00; mem['h7CE2]=8'h00; mem['h7CE3]=8'h00;
    mem['h7CE4]=8'h00; mem['h7CE5]=8'h00; mem['h7CE6]=8'h00; mem['h7CE7]=8'h00;
    mem['h7CE8]=8'h00; mem['h7CE9]=8'h00; mem['h7CEA]=8'h00; mem['h7CEB]=8'h00;
    mem['h7CEC]=8'h00; mem['h7CED]=8'h00; mem['h7CEE]=8'h00; mem['h7CEF]=8'h00;
    mem['h7CF0]=8'h00; mem['h7CF1]=8'h00; mem['h7CF2]=8'h00; mem['h7CF3]=8'h00;
    mem['h7CF4]=8'h00; mem['h7CF5]=8'h00; mem['h7CF6]=8'h00; mem['h7CF7]=8'h00;
    mem['h7CF8]=8'h00; mem['h7CF9]=8'h00; mem['h7CFA]=8'h00; mem['h7CFB]=8'h00;
    mem['h7CFC]=8'h00; mem['h7CFD]=8'h00; mem['h7CFE]=8'h00; mem['h7CFF]=8'h00;
    mem['h7D00]=8'h00; mem['h7D01]=8'h00; mem['h7D02]=8'h00; mem['h7D03]=8'h00;
    mem['h7D04]=8'h00; mem['h7D05]=8'h00; mem['h7D06]=8'h00; mem['h7D07]=8'h00;
    mem['h7D08]=8'h00; mem['h7D09]=8'h00; mem['h7D0A]=8'h00; mem['h7D0B]=8'h00;
    mem['h7D0C]=8'h00; mem['h7D0D]=8'h00; mem['h7D0E]=8'h00; mem['h7D0F]=8'h00;
    mem['h7D10]=8'h00; mem['h7D11]=8'h00; mem['h7D12]=8'h00; mem['h7D13]=8'h00;
    mem['h7D14]=8'h00; mem['h7D15]=8'h00; mem['h7D16]=8'h00; mem['h7D17]=8'h00;
    mem['h7D18]=8'h00; mem['h7D19]=8'h00; mem['h7D1A]=8'h00; mem['h7D1B]=8'h00;
    mem['h7D1C]=8'h00; mem['h7D1D]=8'h00; mem['h7D1E]=8'h00; mem['h7D1F]=8'h00;
    mem['h7D20]=8'h00; mem['h7D21]=8'h00; mem['h7D22]=8'h00; mem['h7D23]=8'h00;
    mem['h7D24]=8'h00; mem['h7D25]=8'h00; mem['h7D26]=8'h00; mem['h7D27]=8'h00;
    mem['h7D28]=8'h00; mem['h7D29]=8'h00; mem['h7D2A]=8'h00; mem['h7D2B]=8'h00;
    mem['h7D2C]=8'h00; mem['h7D2D]=8'h00; mem['h7D2E]=8'h00; mem['h7D2F]=8'h00;
    mem['h7D30]=8'h00; mem['h7D31]=8'h00; mem['h7D32]=8'h00; mem['h7D33]=8'h00;
    mem['h7D34]=8'h00; mem['h7D35]=8'h00; mem['h7D36]=8'h00; mem['h7D37]=8'h00;
    mem['h7D38]=8'h00; mem['h7D39]=8'h00; mem['h7D3A]=8'h00; mem['h7D3B]=8'h00;
    mem['h7D3C]=8'h00; mem['h7D3D]=8'h00; mem['h7D3E]=8'h00; mem['h7D3F]=8'h00;
    mem['h7D40]=8'h00; mem['h7D41]=8'h00; mem['h7D42]=8'h00; mem['h7D43]=8'h00;
    mem['h7D44]=8'h00; mem['h7D45]=8'h00; mem['h7D46]=8'h00; mem['h7D47]=8'h00;
    mem['h7D48]=8'h00; mem['h7D49]=8'h00; mem['h7D4A]=8'h00; mem['h7D4B]=8'h00;
    mem['h7D4C]=8'h00; mem['h7D4D]=8'h00; mem['h7D4E]=8'h00; mem['h7D4F]=8'h00;
    mem['h7D50]=8'h00; mem['h7D51]=8'h00; mem['h7D52]=8'h00; mem['h7D53]=8'h00;
    mem['h7D54]=8'h00; mem['h7D55]=8'h00; mem['h7D56]=8'h00; mem['h7D57]=8'h00;
    mem['h7D58]=8'h00; mem['h7D59]=8'h00; mem['h7D5A]=8'h00; mem['h7D5B]=8'h00;
    mem['h7D5C]=8'h00; mem['h7D5D]=8'h00; mem['h7D5E]=8'h00; mem['h7D5F]=8'h00;
    mem['h7D60]=8'h00; mem['h7D61]=8'h00; mem['h7D62]=8'h00; mem['h7D63]=8'h00;
    mem['h7D64]=8'h00; mem['h7D65]=8'h00; mem['h7D66]=8'h00; mem['h7D67]=8'h00;
    mem['h7D68]=8'h00; mem['h7D69]=8'h00; mem['h7D6A]=8'h00; mem['h7D6B]=8'h00;
    mem['h7D6C]=8'h00; mem['h7D6D]=8'h00; mem['h7D6E]=8'h00; mem['h7D6F]=8'h00;
    mem['h7D70]=8'h00; mem['h7D71]=8'h00; mem['h7D72]=8'h00; mem['h7D73]=8'h00;
    mem['h7D74]=8'h00; mem['h7D75]=8'h00; mem['h7D76]=8'h00; mem['h7D77]=8'h00;
    mem['h7D78]=8'h00; mem['h7D79]=8'h00; mem['h7D7A]=8'h00; mem['h7D7B]=8'h00;
    mem['h7D7C]=8'h00; mem['h7D7D]=8'h00; mem['h7D7E]=8'h00; mem['h7D7F]=8'h00;
    mem['h7D80]=8'h00; mem['h7D81]=8'h00; mem['h7D82]=8'h00; mem['h7D83]=8'h00;
    mem['h7D84]=8'h00; mem['h7D85]=8'h00; mem['h7D86]=8'h00; mem['h7D87]=8'h00;
    mem['h7D88]=8'h00; mem['h7D89]=8'h00; mem['h7D8A]=8'h00; mem['h7D8B]=8'h00;
    mem['h7D8C]=8'h00; mem['h7D8D]=8'h00; mem['h7D8E]=8'h00; mem['h7D8F]=8'h00;
    mem['h7D90]=8'h00; mem['h7D91]=8'h00; mem['h7D92]=8'h00; mem['h7D93]=8'h00;
    mem['h7D94]=8'h00; mem['h7D95]=8'h00; mem['h7D96]=8'h00; mem['h7D97]=8'h00;
    mem['h7D98]=8'h00; mem['h7D99]=8'h00; mem['h7D9A]=8'h00; mem['h7D9B]=8'h00;
    mem['h7D9C]=8'h00; mem['h7D9D]=8'h00; mem['h7D9E]=8'h00; mem['h7D9F]=8'h00;
    mem['h7DA0]=8'h00; mem['h7DA1]=8'h00; mem['h7DA2]=8'h00; mem['h7DA3]=8'h00;
    mem['h7DA4]=8'h00; mem['h7DA5]=8'h00; mem['h7DA6]=8'h00; mem['h7DA7]=8'h00;
    mem['h7DA8]=8'h00; mem['h7DA9]=8'h00; mem['h7DAA]=8'h00; mem['h7DAB]=8'h00;
    mem['h7DAC]=8'h00; mem['h7DAD]=8'h00; mem['h7DAE]=8'h00; mem['h7DAF]=8'h00;
    mem['h7DB0]=8'h00; mem['h7DB1]=8'h00; mem['h7DB2]=8'h00; mem['h7DB3]=8'h00;
    mem['h7DB4]=8'h00; mem['h7DB5]=8'h00; mem['h7DB6]=8'h00; mem['h7DB7]=8'h00;
    mem['h7DB8]=8'h00; mem['h7DB9]=8'h00; mem['h7DBA]=8'h00; mem['h7DBB]=8'h00;
    mem['h7DBC]=8'h00; mem['h7DBD]=8'h00; mem['h7DBE]=8'h00; mem['h7DBF]=8'h00;
    mem['h7DC0]=8'h00; mem['h7DC1]=8'h00; mem['h7DC2]=8'h00; mem['h7DC3]=8'h00;
    mem['h7DC4]=8'h00; mem['h7DC5]=8'h00; mem['h7DC6]=8'h00; mem['h7DC7]=8'h00;
    mem['h7DC8]=8'h00; mem['h7DC9]=8'h00; mem['h7DCA]=8'h00; mem['h7DCB]=8'h00;
    mem['h7DCC]=8'h00; mem['h7DCD]=8'h00; mem['h7DCE]=8'h00; mem['h7DCF]=8'h00;
    mem['h7DD0]=8'h00; mem['h7DD1]=8'h00; mem['h7DD2]=8'h00; mem['h7DD3]=8'h00;
    mem['h7DD4]=8'h00; mem['h7DD5]=8'h00; mem['h7DD6]=8'h00; mem['h7DD7]=8'h00;
    mem['h7DD8]=8'h00; mem['h7DD9]=8'h00; mem['h7DDA]=8'h00; mem['h7DDB]=8'h00;
    mem['h7DDC]=8'h00; mem['h7DDD]=8'h00; mem['h7DDE]=8'h00; mem['h7DDF]=8'h00;
    mem['h7DE0]=8'h00; mem['h7DE1]=8'h00; mem['h7DE2]=8'h00; mem['h7DE3]=8'h00;
    mem['h7DE4]=8'h00; mem['h7DE5]=8'h00; mem['h7DE6]=8'h00; mem['h7DE7]=8'h00;
    mem['h7DE8]=8'h00; mem['h7DE9]=8'h00; mem['h7DEA]=8'h00; mem['h7DEB]=8'h00;
    mem['h7DEC]=8'h00; mem['h7DED]=8'h00; mem['h7DEE]=8'h00; mem['h7DEF]=8'h00;
    mem['h7DF0]=8'h00; mem['h7DF1]=8'h00; mem['h7DF2]=8'h00; mem['h7DF3]=8'h00;
    mem['h7DF4]=8'h00; mem['h7DF5]=8'h00; mem['h7DF6]=8'h00; mem['h7DF7]=8'h00;
    mem['h7DF8]=8'h00; mem['h7DF9]=8'h00; mem['h7DFA]=8'h00; mem['h7DFB]=8'h00;
    mem['h7DFC]=8'h00; mem['h7DFD]=8'h00; mem['h7DFE]=8'h00; mem['h7DFF]=8'h00;
    mem['h7E00]=8'h00; mem['h7E01]=8'h00; mem['h7E02]=8'h00; mem['h7E03]=8'h00;
    mem['h7E04]=8'h00; mem['h7E05]=8'h00; mem['h7E06]=8'h00; mem['h7E07]=8'h00;
    mem['h7E08]=8'h00; mem['h7E09]=8'h00; mem['h7E0A]=8'h00; mem['h7E0B]=8'h00;
    mem['h7E0C]=8'h00; mem['h7E0D]=8'h00; mem['h7E0E]=8'h00; mem['h7E0F]=8'h00;
    mem['h7E10]=8'h00; mem['h7E11]=8'h00; mem['h7E12]=8'h00; mem['h7E13]=8'h00;
    mem['h7E14]=8'h00; mem['h7E15]=8'h00; mem['h7E16]=8'h00; mem['h7E17]=8'h00;
    mem['h7E18]=8'h00; mem['h7E19]=8'h00; mem['h7E1A]=8'h00; mem['h7E1B]=8'h00;
    mem['h7E1C]=8'h00; mem['h7E1D]=8'h00; mem['h7E1E]=8'h00; mem['h7E1F]=8'h00;
    mem['h7E20]=8'h00; mem['h7E21]=8'h00; mem['h7E22]=8'h00; mem['h7E23]=8'h00;
    mem['h7E24]=8'h00; mem['h7E25]=8'h00; mem['h7E26]=8'h00; mem['h7E27]=8'h00;
    mem['h7E28]=8'h00; mem['h7E29]=8'h00; mem['h7E2A]=8'h00; mem['h7E2B]=8'h00;
    mem['h7E2C]=8'h00; mem['h7E2D]=8'h00; mem['h7E2E]=8'h00; mem['h7E2F]=8'h00;
    mem['h7E30]=8'h00; mem['h7E31]=8'h00; mem['h7E32]=8'h00; mem['h7E33]=8'h00;
    mem['h7E34]=8'h00; mem['h7E35]=8'h00; mem['h7E36]=8'h00; mem['h7E37]=8'h00;
    mem['h7E38]=8'h00; mem['h7E39]=8'h00; mem['h7E3A]=8'h00; mem['h7E3B]=8'h00;
    mem['h7E3C]=8'h00; mem['h7E3D]=8'h00; mem['h7E3E]=8'h00; mem['h7E3F]=8'h00;
    mem['h7E40]=8'h00; mem['h7E41]=8'h00; mem['h7E42]=8'h00; mem['h7E43]=8'h00;
    mem['h7E44]=8'h00; mem['h7E45]=8'h00; mem['h7E46]=8'h00; mem['h7E47]=8'h00;
    mem['h7E48]=8'h00; mem['h7E49]=8'h00; mem['h7E4A]=8'h00; mem['h7E4B]=8'h00;
    mem['h7E4C]=8'h00; mem['h7E4D]=8'h00; mem['h7E4E]=8'h00; mem['h7E4F]=8'h00;
    mem['h7E50]=8'h00; mem['h7E51]=8'h00; mem['h7E52]=8'h00; mem['h7E53]=8'h00;
    mem['h7E54]=8'h00; mem['h7E55]=8'h00; mem['h7E56]=8'h00; mem['h7E57]=8'h00;
    mem['h7E58]=8'h00; mem['h7E59]=8'h00; mem['h7E5A]=8'h00; mem['h7E5B]=8'h00;
    mem['h7E5C]=8'h00; mem['h7E5D]=8'h00; mem['h7E5E]=8'h00; mem['h7E5F]=8'h00;
    mem['h7E60]=8'h00; mem['h7E61]=8'h00; mem['h7E62]=8'h00; mem['h7E63]=8'h00;
    mem['h7E64]=8'h00; mem['h7E65]=8'h00; mem['h7E66]=8'h00; mem['h7E67]=8'h00;
    mem['h7E68]=8'h00; mem['h7E69]=8'h00; mem['h7E6A]=8'h00; mem['h7E6B]=8'h00;
    mem['h7E6C]=8'h00; mem['h7E6D]=8'h00; mem['h7E6E]=8'h00; mem['h7E6F]=8'h00;
    mem['h7E70]=8'h00; mem['h7E71]=8'h00; mem['h7E72]=8'h00; mem['h7E73]=8'h00;
    mem['h7E74]=8'h00; mem['h7E75]=8'h00; mem['h7E76]=8'h00; mem['h7E77]=8'h00;
    mem['h7E78]=8'h00; mem['h7E79]=8'h00; mem['h7E7A]=8'h00; mem['h7E7B]=8'h00;
    mem['h7E7C]=8'h00; mem['h7E7D]=8'h00; mem['h7E7E]=8'h00; mem['h7E7F]=8'h00;
    mem['h7E80]=8'h00; mem['h7E81]=8'h00; mem['h7E82]=8'h00; mem['h7E83]=8'h00;
    mem['h7E84]=8'h00; mem['h7E85]=8'h00; mem['h7E86]=8'h00; mem['h7E87]=8'h00;
    mem['h7E88]=8'h00; mem['h7E89]=8'h00; mem['h7E8A]=8'h00; mem['h7E8B]=8'h00;
    mem['h7E8C]=8'h00; mem['h7E8D]=8'h00; mem['h7E8E]=8'h00; mem['h7E8F]=8'h00;
    mem['h7E90]=8'h00; mem['h7E91]=8'h00; mem['h7E92]=8'h00; mem['h7E93]=8'h00;
    mem['h7E94]=8'h00; mem['h7E95]=8'h00; mem['h7E96]=8'h00; mem['h7E97]=8'h00;
    mem['h7E98]=8'h00; mem['h7E99]=8'h00; mem['h7E9A]=8'h00; mem['h7E9B]=8'h00;
    mem['h7E9C]=8'h00; mem['h7E9D]=8'h00; mem['h7E9E]=8'h00; mem['h7E9F]=8'h00;
    mem['h7EA0]=8'h00; mem['h7EA1]=8'h00; mem['h7EA2]=8'h00; mem['h7EA3]=8'h00;
    mem['h7EA4]=8'h00; mem['h7EA5]=8'h00; mem['h7EA6]=8'h00; mem['h7EA7]=8'h00;
    mem['h7EA8]=8'h00; mem['h7EA9]=8'h00; mem['h7EAA]=8'h00; mem['h7EAB]=8'h00;
    mem['h7EAC]=8'h00; mem['h7EAD]=8'h00; mem['h7EAE]=8'h00; mem['h7EAF]=8'h00;
    mem['h7EB0]=8'h00; mem['h7EB1]=8'h00; mem['h7EB2]=8'h00; mem['h7EB3]=8'h00;
    mem['h7EB4]=8'h00; mem['h7EB5]=8'h00; mem['h7EB6]=8'h00; mem['h7EB7]=8'h00;
    mem['h7EB8]=8'h00; mem['h7EB9]=8'h00; mem['h7EBA]=8'h00; mem['h7EBB]=8'h00;
    mem['h7EBC]=8'h00; mem['h7EBD]=8'h00; mem['h7EBE]=8'h00; mem['h7EBF]=8'h00;
    mem['h7EC0]=8'h00; mem['h7EC1]=8'h00; mem['h7EC2]=8'h00; mem['h7EC3]=8'h00;
    mem['h7EC4]=8'h00; mem['h7EC5]=8'h00; mem['h7EC6]=8'h00; mem['h7EC7]=8'h00;
    mem['h7EC8]=8'h00; mem['h7EC9]=8'h00; mem['h7ECA]=8'h00; mem['h7ECB]=8'h00;
    mem['h7ECC]=8'h00; mem['h7ECD]=8'h00; mem['h7ECE]=8'h00; mem['h7ECF]=8'h00;
    mem['h7ED0]=8'h00; mem['h7ED1]=8'h00; mem['h7ED2]=8'h00; mem['h7ED3]=8'h00;
    mem['h7ED4]=8'h00; mem['h7ED5]=8'h00; mem['h7ED6]=8'h00; mem['h7ED7]=8'h00;
    mem['h7ED8]=8'h00; mem['h7ED9]=8'h00; mem['h7EDA]=8'h00; mem['h7EDB]=8'h00;
    mem['h7EDC]=8'h00; mem['h7EDD]=8'h00; mem['h7EDE]=8'h00; mem['h7EDF]=8'h00;
    mem['h7EE0]=8'h00; mem['h7EE1]=8'h00; mem['h7EE2]=8'h00; mem['h7EE3]=8'h00;
    mem['h7EE4]=8'h00; mem['h7EE5]=8'h00; mem['h7EE6]=8'h00; mem['h7EE7]=8'h00;
    mem['h7EE8]=8'h00; mem['h7EE9]=8'h00; mem['h7EEA]=8'h00; mem['h7EEB]=8'h00;
    mem['h7EEC]=8'h00; mem['h7EED]=8'h00; mem['h7EEE]=8'h00; mem['h7EEF]=8'h00;
    mem['h7EF0]=8'h00; mem['h7EF1]=8'h00; mem['h7EF2]=8'h00; mem['h7EF3]=8'h00;
    mem['h7EF4]=8'h00; mem['h7EF5]=8'h00; mem['h7EF6]=8'h00; mem['h7EF7]=8'h00;
    mem['h7EF8]=8'h00; mem['h7EF9]=8'h00; mem['h7EFA]=8'h00; mem['h7EFB]=8'h00;
    mem['h7EFC]=8'h00; mem['h7EFD]=8'h00; mem['h7EFE]=8'h00; mem['h7EFF]=8'h00;
    mem['h7F00]=8'h00; mem['h7F01]=8'h00; mem['h7F02]=8'h00; mem['h7F03]=8'h00;
    mem['h7F04]=8'h00; mem['h7F05]=8'h00; mem['h7F06]=8'h00; mem['h7F07]=8'h00;
    mem['h7F08]=8'h00; mem['h7F09]=8'h00; mem['h7F0A]=8'h00; mem['h7F0B]=8'h00;
    mem['h7F0C]=8'h00; mem['h7F0D]=8'h00; mem['h7F0E]=8'h00; mem['h7F0F]=8'h00;
    mem['h7F10]=8'h00; mem['h7F11]=8'h00; mem['h7F12]=8'h00; mem['h7F13]=8'h00;
    mem['h7F14]=8'h00; mem['h7F15]=8'h00; mem['h7F16]=8'h00; mem['h7F17]=8'h00;
    mem['h7F18]=8'h00; mem['h7F19]=8'h00; mem['h7F1A]=8'h00; mem['h7F1B]=8'h00;
    mem['h7F1C]=8'h00; mem['h7F1D]=8'h00; mem['h7F1E]=8'h00; mem['h7F1F]=8'h00;
    mem['h7F20]=8'h00; mem['h7F21]=8'h00; mem['h7F22]=8'h00; mem['h7F23]=8'h00;
    mem['h7F24]=8'h00; mem['h7F25]=8'h00; mem['h7F26]=8'h00; mem['h7F27]=8'h00;
    mem['h7F28]=8'h00; mem['h7F29]=8'h00; mem['h7F2A]=8'h00; mem['h7F2B]=8'h00;
    mem['h7F2C]=8'h00; mem['h7F2D]=8'h00; mem['h7F2E]=8'h00; mem['h7F2F]=8'h00;
    mem['h7F30]=8'h00; mem['h7F31]=8'h00; mem['h7F32]=8'h00; mem['h7F33]=8'h00;
    mem['h7F34]=8'h00; mem['h7F35]=8'h00; mem['h7F36]=8'h00; mem['h7F37]=8'h00;
    mem['h7F38]=8'h00; mem['h7F39]=8'h00; mem['h7F3A]=8'h00; mem['h7F3B]=8'h00;
    mem['h7F3C]=8'h00; mem['h7F3D]=8'h00; mem['h7F3E]=8'h00; mem['h7F3F]=8'h00;
    mem['h7F40]=8'h00; mem['h7F41]=8'h00; mem['h7F42]=8'h00; mem['h7F43]=8'h00;
    mem['h7F44]=8'h00; mem['h7F45]=8'h00; mem['h7F46]=8'h00; mem['h7F47]=8'h00;
    mem['h7F48]=8'h00; mem['h7F49]=8'h00; mem['h7F4A]=8'h00; mem['h7F4B]=8'h00;
    mem['h7F4C]=8'h00; mem['h7F4D]=8'h00; mem['h7F4E]=8'h00; mem['h7F4F]=8'h00;
    mem['h7F50]=8'h00; mem['h7F51]=8'h00; mem['h7F52]=8'h00; mem['h7F53]=8'h00;
    mem['h7F54]=8'h00; mem['h7F55]=8'h00; mem['h7F56]=8'h00; mem['h7F57]=8'h00;
    mem['h7F58]=8'h00; mem['h7F59]=8'h00; mem['h7F5A]=8'h00; mem['h7F5B]=8'h00;
    mem['h7F5C]=8'h00; mem['h7F5D]=8'h00; mem['h7F5E]=8'h00; mem['h7F5F]=8'h00;
    mem['h7F60]=8'h00; mem['h7F61]=8'h00; mem['h7F62]=8'h00; mem['h7F63]=8'h00;
    mem['h7F64]=8'h00; mem['h7F65]=8'h00; mem['h7F66]=8'h00; mem['h7F67]=8'h00;
    mem['h7F68]=8'h00; mem['h7F69]=8'h00; mem['h7F6A]=8'h00; mem['h7F6B]=8'h00;
    mem['h7F6C]=8'h00; mem['h7F6D]=8'h00; mem['h7F6E]=8'h00; mem['h7F6F]=8'h00;
    mem['h7F70]=8'h00; mem['h7F71]=8'h00; mem['h7F72]=8'h00; mem['h7F73]=8'h00;
    mem['h7F74]=8'h00; mem['h7F75]=8'h00; mem['h7F76]=8'h00; mem['h7F77]=8'h00;
    mem['h7F78]=8'h00; mem['h7F79]=8'h00; mem['h7F7A]=8'h00; mem['h7F7B]=8'h00;
    mem['h7F7C]=8'h00; mem['h7F7D]=8'h00; mem['h7F7E]=8'h00; mem['h7F7F]=8'h00;
    mem['h7F80]=8'h00; mem['h7F81]=8'h00; mem['h7F82]=8'h00; mem['h7F83]=8'h00;
    mem['h7F84]=8'h00; mem['h7F85]=8'h00; mem['h7F86]=8'h00; mem['h7F87]=8'h00;
    mem['h7F88]=8'h00; mem['h7F89]=8'h00; mem['h7F8A]=8'h00; mem['h7F8B]=8'h00;
    mem['h7F8C]=8'h00; mem['h7F8D]=8'h00; mem['h7F8E]=8'h00; mem['h7F8F]=8'h00;
    mem['h7F90]=8'h00; mem['h7F91]=8'h00; mem['h7F92]=8'h00; mem['h7F93]=8'h00;
    mem['h7F94]=8'h00; mem['h7F95]=8'h00; mem['h7F96]=8'h00; mem['h7F97]=8'h00;
    mem['h7F98]=8'h00; mem['h7F99]=8'h00; mem['h7F9A]=8'h00; mem['h7F9B]=8'h00;
    mem['h7F9C]=8'h00; mem['h7F9D]=8'h00; mem['h7F9E]=8'h00; mem['h7F9F]=8'h00;
    mem['h7FA0]=8'h00; mem['h7FA1]=8'h00; mem['h7FA2]=8'h00; mem['h7FA3]=8'h00;
    mem['h7FA4]=8'h00; mem['h7FA5]=8'h00; mem['h7FA6]=8'h00; mem['h7FA7]=8'h00;
    mem['h7FA8]=8'h00; mem['h7FA9]=8'h00; mem['h7FAA]=8'h00; mem['h7FAB]=8'h00;
    mem['h7FAC]=8'h00; mem['h7FAD]=8'h00; mem['h7FAE]=8'h00; mem['h7FAF]=8'h00;
    mem['h7FB0]=8'h00; mem['h7FB1]=8'h00; mem['h7FB2]=8'h00; mem['h7FB3]=8'h00;
    mem['h7FB4]=8'h00; mem['h7FB5]=8'h00; mem['h7FB6]=8'h00; mem['h7FB7]=8'h00;
    mem['h7FB8]=8'h00; mem['h7FB9]=8'h00; mem['h7FBA]=8'h00; mem['h7FBB]=8'h00;
    mem['h7FBC]=8'h00; mem['h7FBD]=8'h00; mem['h7FBE]=8'h00; mem['h7FBF]=8'h00;
    mem['h7FC0]=8'h00; mem['h7FC1]=8'h00; mem['h7FC2]=8'h00; mem['h7FC3]=8'h00;
    mem['h7FC4]=8'h00; mem['h7FC5]=8'h00; mem['h7FC6]=8'h00; mem['h7FC7]=8'h00;
    mem['h7FC8]=8'h00; mem['h7FC9]=8'h00; mem['h7FCA]=8'h00; mem['h7FCB]=8'h00;
    mem['h7FCC]=8'h00; mem['h7FCD]=8'h00; mem['h7FCE]=8'h00; mem['h7FCF]=8'h00;
    mem['h7FD0]=8'h00; mem['h7FD1]=8'h00; mem['h7FD2]=8'h00; mem['h7FD3]=8'h00;
    mem['h7FD4]=8'h00; mem['h7FD5]=8'h00; mem['h7FD6]=8'h00; mem['h7FD7]=8'h00;
    mem['h7FD8]=8'h00; mem['h7FD9]=8'h00; mem['h7FDA]=8'h00; mem['h7FDB]=8'h00;
    mem['h7FDC]=8'h00; mem['h7FDD]=8'h00; mem['h7FDE]=8'h00; mem['h7FDF]=8'h00;
    mem['h7FE0]=8'h00; mem['h7FE1]=8'h00; mem['h7FE2]=8'h00; mem['h7FE3]=8'h00;
    mem['h7FE4]=8'h00; mem['h7FE5]=8'h00; mem['h7FE6]=8'h00; mem['h7FE7]=8'h00;
    mem['h7FE8]=8'h00; mem['h7FE9]=8'h00; mem['h7FEA]=8'h00; mem['h7FEB]=8'h00;
    mem['h7FEC]=8'h00; mem['h7FED]=8'h00; mem['h7FEE]=8'h00; mem['h7FEF]=8'h00;
    mem['h7FF0]=8'h00; mem['h7FF1]=8'h00; mem['h7FF2]=8'h00; mem['h7FF3]=8'h00;
    mem['h7FF4]=8'h00; mem['h7FF5]=8'h00; mem['h7FF6]=8'h00; mem['h7FF7]=8'h00;
    mem['h7FF8]=8'h00; mem['h7FF9]=8'h00; mem['h7FFA]=8'h00; mem['h7FFB]=8'h00;
    mem['h7FFC]=8'h00; mem['h7FFD]=8'h00; mem['h7FFE]=8'h00; mem['h7FFF]=8'h00;
end
